--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : ssm_demo.vh
--FILE GENERATED ON : Fri Mar 12 09:18:02 2010

a2rtap.vhd
cmpr.vhd
dsp.vhd
dummy_unit_synth_removes.vhd
eu.vhd
h264.vhd
host_processor.vhd
im.vhd
mcb.vhd
me.vhd
pc.vhd
rf.vhd
ssm_demo.vhd
ssm_master.vhd
wb.vhd
