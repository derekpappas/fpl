`include "defines.v"

module u1();
// Location of source csl unit: file name = ar16.csl line number = 35
  `include "u1.logic.v"
endmodule

