// Test type: net_assignment - binary operator, 1 attribute instance
// Vparser rule name:
// Author: andreib
module netasign6;
wire a,b,c,d;
assign a=b*(*c*)d;
endmodule
