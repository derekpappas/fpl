`ifndef DFF_NS
`define DFF_NS

module dff_ns;
endmodule

module dffrl_async_ns;
endmodule

module dffrle_ns;
endmodule

module dffrl_ns;
endmodule

module dffsl_async_ns;
endmodule

module ucb_bus_out;
endmodule

module ucb_bus_in;
endmodule

`endif
