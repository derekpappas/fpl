//test type : specify_block_declaration
//author : Dramba Doru-Gabriel
module specify_block_data_event0(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event2(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event3(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event4(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event5(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event6(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event7(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event8(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event9(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event10(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event11(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event12(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event13(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event14(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event15(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event16(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event17(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event18(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event19(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event20(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event21(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event22(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event23(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event24(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event25(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event26(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event27(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event28(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event29(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event30(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event31(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event32(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event33(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event34(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event35(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event36(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event37(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event38(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event39(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event40(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event41(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event42(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event43(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event44(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event45(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event46(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event47(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event48(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event49(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event50(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event51(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event52(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event53(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event54(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event55(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event56(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event57(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event58(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event59(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event60(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event61(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event62(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event63(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event64(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event65(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event66(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event67(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event68(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event69(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event70(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event71(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event72(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event73(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event74(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event75(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event76(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event77(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event78(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event79(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event80(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event81(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event82(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event83(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event84(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event85(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event86(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event87(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event88(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event89(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event90(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event91(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event92(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event93(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event94(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event95(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event96(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event97(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event98(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event99(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event100(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event101(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event102(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event103(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event104(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event105(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event106(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event107(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event108(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event109(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event110(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event111(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event112(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event113(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event114(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event115(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event116(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event117(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event118(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event119(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event120(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event121(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event122(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event123(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event124(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event125(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event126(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event127(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event128(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event129(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event130(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event131(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event132(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event133(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event134(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event135(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event136(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event137(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event138(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event139(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event140(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event141(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event142(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event143(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event144(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event145(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event146(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event147(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event148(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event149(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event150(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event151(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event152(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event153(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event154(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event155(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event156(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event157(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event158(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event159(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event160(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event161(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event162(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event163(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event164(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event165(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event166(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event167(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event168(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event169(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event170(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event171(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event172(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event173(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event174(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event175(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event176(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event177(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event178(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event179(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event180(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event181(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event182(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event183(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event184(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event185(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event186(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event187(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event188(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event189(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event190(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event191(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event192(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event193(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event194(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event195(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event196(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event197(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event198(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event199(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event200(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event201(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event202(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event203(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event204(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event205(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event206(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event207(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event208(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event209(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event210(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event211(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event212(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event213(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event214(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event215(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event216(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event217(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event218(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event219(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event220(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event221(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event222(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event223(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event224(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event225(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event226(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event227(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event228(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event229(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event230(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event231(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event232(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event233(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event234(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event235(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event236(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event237(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event238(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event239(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event240(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event241(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event242(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event243(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event244(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event245(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event246(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event247(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event248(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event249(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event250(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event251(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event252(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event253(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event254(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event255(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event256(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event257(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event258(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event259(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event260(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event261(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event262(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event263(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event264(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event265(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event266(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event267(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event268(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event269(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event270(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event271(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event272(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event273(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event274(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event275(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event276(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event277(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event278(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event279(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event280(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event281(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event282(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event283(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event284(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event285(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event286(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event287(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event288(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event289(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event290(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event291(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event292(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event293(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event294(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event295(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event296(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event297(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event298(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event299(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event300(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event301(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event302(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event303(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event304(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event305(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event306(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event307(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event308(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event309(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event310(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event311(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( posedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event312(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event313(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event314(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event315(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event316(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event317(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event318(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event319(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event320(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event321(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event322(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event323(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event324(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event325(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event326(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event327(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event328(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event329(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event330(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event331(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event332(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event333(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event334(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event335(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event336(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event337(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event338(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event339(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event340(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event341(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event342(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event343(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event344(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event345(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event346(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event347(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event348(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event349(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event350(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event351(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event352(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event353(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event354(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event355(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event356(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event357(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event358(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event359(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event360(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event361(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event362(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event363(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event364(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event365(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event366(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event367(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event368(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event369(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event370(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event371(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event372(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event373(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event374(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event375(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event376(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event377(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event378(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event379(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event380(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event381(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event382(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event383(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event384(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event385(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event386(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event387(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event388(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event389(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event390(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event391(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event392(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event393(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event394(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event395(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event396(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event397(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event398(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event399(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event400(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event401(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event402(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event403(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event404(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event405(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event406(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event407(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event408(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event409(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event410(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event411(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event412(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event413(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event414(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event415(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event416(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event417(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event418(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event419(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event420(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event421(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event422(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event423(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event424(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event425(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event426(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event427(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event428(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event429(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event430(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event431(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event432(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event433(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event434(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event435(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event436(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event437(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event438(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event439(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event440(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event441(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event442(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event443(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event444(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event445(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event446(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event447(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event448(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event449(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event450(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event451(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event452(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event453(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event454(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event455(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event456(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event457(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event458(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event459(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event460(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event461(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event462(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event463(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event464(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event465(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event466(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event467(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( negedge inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event468(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event469(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event470(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event471(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event472(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event473(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event474(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event475(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event476(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event477(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event478(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event479(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event480(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event481(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event482(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event483(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event484(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event485(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event486(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event487(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event488(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event489(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event490(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event491(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event492(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event493(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event494(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event495(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event496(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event497(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event498(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event499(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event500(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event501(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event502(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event503(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event504(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event505(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event506(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event507(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event508(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event509(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event510(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event511(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event512(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event513(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event514(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event515(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event516(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event517(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event518(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event519(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event520(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event521(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event522(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event523(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event524(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event525(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event526(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event527(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event528(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event529(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event530(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event531(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event532(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event533(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event534(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event535(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event536(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event537(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event538(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event539(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event540(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event541(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event542(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event543(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event544(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event545(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event546(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event547(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event548(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event549(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event550(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event551(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event552(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event553(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event554(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event555(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event556(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event557(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event558(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event559(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event560(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event561(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event562(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event563(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event564(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event565(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event566(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event567(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event568(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event569(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event570(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event571(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event572(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event573(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event574(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event575(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event576(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event577(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event578(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event579(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event580(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event581(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event582(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event583(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event584(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event585(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event586(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event587(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event588(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event589(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event590(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event591(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event592(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event593(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event594(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event595(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event596(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event597(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event598(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event599(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event600(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event601(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event602(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event603(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event604(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event605(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event606(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event607(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event608(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event609(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event610(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event611(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event612(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event613(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event614(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event615(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event616(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event617(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event618(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event619(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event620(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event621(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event622(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event623(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 01 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event624(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event625(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event626(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event627(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event628(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event629(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event630(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event631(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event632(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event633(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event634(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event635(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event636(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event637(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event638(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event639(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event640(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event641(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event642(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event643(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event644(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event645(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event646(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event647(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event648(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event649(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event650(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event651(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event652(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event653(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event654(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event655(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event656(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event657(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event658(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event659(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event660(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event661(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event662(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event663(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event664(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event665(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event666(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event667(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event668(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event669(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event670(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event671(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event672(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event673(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event674(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event675(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event676(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event677(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event678(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event679(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event680(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event681(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event682(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event683(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event684(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event685(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event686(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event687(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event688(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event689(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event690(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event691(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event692(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event693(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event694(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event695(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event696(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event697(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event698(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event699(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event700(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event701(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event702(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event703(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event704(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event705(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event706(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event707(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event708(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event709(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event710(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event711(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event712(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event713(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event714(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event715(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event716(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event717(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event718(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event719(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event720(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event721(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event722(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event723(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event724(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event725(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event726(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event727(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event728(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event729(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event730(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event731(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event732(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event733(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event734(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event735(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event736(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event737(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event738(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event739(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event740(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event741(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event742(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event743(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event744(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event745(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event746(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event747(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event748(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event749(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event750(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event751(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event752(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event753(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event754(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event755(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event756(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event757(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event758(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event759(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event760(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event761(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event762(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event763(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event764(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event765(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event766(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event767(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event768(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event769(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event770(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event771(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event772(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event773(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event774(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event775(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event776(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event777(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event778(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event779(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 10 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event780(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event781(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event782(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event783(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event784(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event785(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event786(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event787(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event788(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event789(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event790(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event791(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event792(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event793(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event794(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event795(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event796(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event797(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event798(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event799(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event800(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event801(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event802(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event803(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event804(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event805(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event806(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event807(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event808(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event809(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event810(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event811(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event812(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event813(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event814(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event815(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event816(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event817(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event818(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event819(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event820(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event821(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event822(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event823(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event824(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event825(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event826(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event827(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event828(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event829(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event830(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event831(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event832(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event833(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event834(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event835(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event836(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event837(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event838(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event839(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event840(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event841(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event842(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event843(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event844(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event845(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event846(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event847(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event848(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event849(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event850(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event851(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event852(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event853(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event854(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event855(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event856(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event857(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event858(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event859(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event860(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event861(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event862(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event863(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event864(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event865(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event866(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event867(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event868(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event869(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event870(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event871(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event872(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event873(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event874(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event875(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event876(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event877(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event878(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event879(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event880(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event881(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event882(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event883(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event884(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event885(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event886(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event887(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event888(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event889(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event890(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event891(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event892(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event893(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event894(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event895(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event896(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event897(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event898(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event899(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event900(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event901(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event902(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event903(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event904(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event905(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event906(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event907(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event908(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event909(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event910(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event911(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event912(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event913(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event914(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event915(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event916(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event917(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event918(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event919(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event920(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event921(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event922(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event923(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event924(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event925(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event926(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event927(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event928(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event929(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event930(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event931(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event932(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event933(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event934(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event935(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ 0X ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event936(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event937(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event938(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event939(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event940(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event941(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event942(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event943(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event944(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event945(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event946(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event947(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event948(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event949(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event950(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event951(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event952(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event953(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event954(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event955(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event956(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event957(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event958(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event959(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event960(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event961(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event962(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event963(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event964(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event965(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event966(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event967(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event968(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event969(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event970(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event971(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event972(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event973(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event974(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event975(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event976(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event977(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event978(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event979(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event980(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event981(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event982(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event983(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event984(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event985(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event986(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event987(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event988(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event989(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event990(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event991(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event992(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event993(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event994(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event995(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event996(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event997(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event998(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event999(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1000(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1001(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1002(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1003(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1004(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1005(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1006(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1007(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1008(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1009(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1010(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1011(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1012(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1013(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1014(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1015(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1016(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1017(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1018(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1019(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1020(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1021(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1022(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1023(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1024(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1025(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1026(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1027(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1028(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1029(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1030(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1031(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1032(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1033(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1034(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1035(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1036(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1037(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1038(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1039(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1040(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1041(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1042(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1043(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1044(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1045(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1046(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1047(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1048(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1049(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1050(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1051(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1052(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1053(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1054(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1055(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1056(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1057(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1058(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1059(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1060(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1061(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1062(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1063(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1064(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1065(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1066(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1067(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1068(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1069(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1070(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1071(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1072(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1073(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1074(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1075(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1076(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1077(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1078(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1079(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1080(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1081(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1082(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1083(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1084(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1085(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1086(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1087(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1088(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1089(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1090(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1091(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ x0 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1092(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1093(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1094(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1095(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1096(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1097(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1098(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1099(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1100(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1101(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1102(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1103(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1104(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1105(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1106(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1107(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1108(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1109(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1110(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1111(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1112(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1113(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1114(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1115(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1116(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1117(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1118(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1119(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1120(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1121(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1122(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1123(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1124(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1125(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1126(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1127(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ~exp , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1128(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1129(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1130(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1131(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1132(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1133(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1134(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1135(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1136(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1137(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1138(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1139(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp==1'b0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1140(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1141(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1142(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1143(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1144(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1145(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1146(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1147(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1148(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1149(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1150(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1151(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp===1'b1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1152(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1153(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1154(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1155(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1156(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1157(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1158(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1159(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1160(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1161(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1162(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1163(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!='B0 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1164(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1165(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1166(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1167(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1168(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1169(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1170(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1171(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1172(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1173(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1174(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1175(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& exp!=='B1 , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1176(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1177(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1178(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1179(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1180(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1181(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1182(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1183(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1184(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1185(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1186(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1187(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1188(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1189(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1190(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1191(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1192(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1193(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1194(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1195(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1196(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1197(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1198(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1199(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( ~exp ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1200(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1201(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1202(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1203(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1204(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1205(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1206(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1207(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1208(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1209(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1210(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1211(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp==1'b0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1212(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1213(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1214(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1215(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1216(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1217(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1218(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1219(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1220(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1221(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1222(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1223(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp===1'b1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1224(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1225(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1226(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1227(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1228(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1229(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1230(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1231(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1232(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1233(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1234(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1235(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!='B0 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1236(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1237(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1238(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1239(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1240(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1241(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1242(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1243(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1244(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier , "timing_check_limit" , notify_reg ); endspecify
endmodule
module specify_block_data_event1245(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" ); endspecify
endmodule
module specify_block_data_event1246(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , ); endspecify
endmodule
module specify_block_data_event1247(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setup( edge[ Z1 ] inoutPortIdentifier &&& ( exp!=='B1 ) , posedge inoutPortIdentifier &&& exp , "timing_check_limit" , notify_reg ); endspecify
endmodule
