-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_mbist_cslc_generated/code/vhdl/u_alu.vhd
-- FILE GENERATED ON : Tue Feb 17 20:24:21 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_alu\ is
  port(\p_op1\ : in csl_bit_vector(10#15# downto 10#0#);
       \p_op2\ : in csl_bit_vector(10#15# downto 10#0#);
       \p_opsel\ : in csl_bit_vector(10#2# downto 10#0#);
       \p_cin\ : in csl_bit;
       \p_res\ : out csl_bit_vector(10#15# downto 10#0#);
       \p_cout\ : out csl_bit);
begin
end entity;

architecture \u_alu_logic\ of \u_alu\ is
begin
end architecture;

