-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top_cslc_generated/code/vhdl/c.vhd
-- FILE GENERATED ON : Mon Feb 16 21:21:57 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \c\ is
  port(\c_in\ : in csl_bit;
       \c_out\ : out csl_bit_vector(10#16# - 10#1# downto 10#0#));
begin
end entity;

architecture \c_logic\ of \c\ is
begin
end architecture;

