//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2005, 2006, 2007 FastpathLogic Inc

module u();
  wire sgg0_sg0_s1;
  wire sgg0_sg0_s2;
  wire sgg0_sg0_s3;
  wire sgg0_s4;
endmodule

