// Test type: par_block - fork - join
// Vparser rule name:
// Author: andreib
module par_block1;
initial fork join
endmodule
