`include "defines.v"

module l0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 79
  input [1 - 1:0] ar_sa0_s10;
  k0 k0(.ar_sa0_s10(ar_sa0_s10));
  `include "l0.logic.vh"
endmodule

