//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : u.v
//FILE GENERATED ON : Fri Oct 26 14:45:17 2007

module u(p1,
         p2,
         p3);
// Location of source csl unit: file name =  line number = 1
  input p1;
  input p2;
  output p3;
endmodule

