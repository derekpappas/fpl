proc.vhd
cluster.vhd
