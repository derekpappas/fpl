// Test type: Real numbers - underscores within
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1234567.12e1_23_;
endmodule
