//test type : {module_path_expression}
//vparser rule name : 
//author : Bogdan Mereghea
module module_path_concatenation1;
    wire a;
    assign a = {{1'b1}};
endmodule
