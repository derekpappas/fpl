`include "defines.v"

module i0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 55
  input [1 - 1:0] ar_sa0_s10;
  h0 h0(.ar_sa0_s10(ar_sa0_s10));
  `include "i0.logic.vh"
endmodule

