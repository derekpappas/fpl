module a(x);
output reg x = 1'b1;
endmodule 

module b(x);
input x;
endmodule