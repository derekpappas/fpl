//test type : non_port_module_item ::= local_parameter_declaration
//vparser rule name : 
//author : Codrin
module test_0370;
 (* debug = 0, test, sign *)
 localparam size = 7;
endmodule
