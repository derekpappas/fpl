//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : ddr_buf_ctrl.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module ddr_buf_ctrl(lbdummy2,
                    dc_dbcdummy5);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 11
  input lbdummy2;
  input dc_dbcdummy5;
  `include "ddr_buf_ctrl.logic.v"
endmodule

