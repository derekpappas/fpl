//test type : module_declaration
//vparser rule name : 
//author : Codrin
(* a *)
(* a = 1 *)
(* a, b *)
(* a = 1, b *)
(* a, b = 1 *)
(* a = 1, b = 1 *)
(* a, b, c *)
module declaration_060;
endmodule
