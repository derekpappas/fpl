// Test type: procedural continuous assignment - force variable assignment
// Vparser rule name:
// Author: andreib
module procedural_continuous_assignment3;
reg a;
initial force a=1;
endmodule
