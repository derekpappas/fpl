//test type : module_or_generate_item ::= module_or_generate_item_declaration (net_declaration)
//vparser rule name : 
//author : Codrin
module test_0170;
 (* nets = 1 *) wire [7:0] out;
endmodule
