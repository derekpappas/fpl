mem.vhd
u.vhd
