`include "defines.v"

module pc();
// Location of source csl unit: file name = /Volumes/s2/unfuddle_ssm_repo/ssm_ssmrepo/ssm/hw/ssm/ssm_demo.csl line number = 95
  `include "pc.logic.vh"
endmodule

