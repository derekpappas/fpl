module prefix();
    parameter WIDTH=4;
    parameter DEPTH=8;
    
    ETICHETA 
    reg [WIDTH-1:0] as[0:DEPTH-1];
endmodule