`include "defines.v"

module v0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 150
  input [1 - 1:0] ar_sa0_s10;
  u0 u0(.ar_sa0_s10(ar_sa0_s10));
  `include "v0.logic.vh"
endmodule

