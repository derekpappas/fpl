// Test type: par_block - fork - block.id (ASCII) - join
// Vparser rule name:
// Author: andreib
module par_block2;
initial fork:abcdefghijklmnopqrstuvwxyzABCDEFGHIJKLMNOPQRSTUVWXYZ1234567890_$ join
endmodule
