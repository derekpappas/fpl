// Test type: seq_block - begin - block.id (ASCII) - end
// Vparser rule name:
// Author: andreib
module seq_block2;
initial begin:abcdefghijklmnopqrstuvwxyzABCDEFGHIJKLMNOPQRSTUVWXYZ1234567890_$ end
endmodule
