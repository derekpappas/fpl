`include "defines.v"

module s1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 292
  output [1 - 1:0] ar_sa0_s10;
  r1 r10(.ar_sa0_s10(ar_sa0_s10));
  `include "s1.logic.vh"
endmodule

