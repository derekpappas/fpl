module u1();
    u1 u11();
    u2 u2();
endmodule

module u2();
endmodule