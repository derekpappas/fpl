//test type : module_or_generate_item ::= operator
//vparser rule name : 
//author : Codrin
module test_0300(input c, output a);
 wire b;
 assign a = b + (* xmodel ="cla" *) c;
endmodule
