-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top_cslc_generated/code/vhdl/u_c.vhd
-- FILE GENERATED ON : Wed Mar 11 20:22:38 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_c\ is
  port(\ck\ : in csl_bit;
       \reset\ : in csl_bit;
       \p_c_in\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \p_c_out\ : out csl_bit_vector(10#8# - 10#1# downto 10#0#));
begin
end entity;

architecture \u_c_logic\ of \u_c\ is
begin
end architecture;

