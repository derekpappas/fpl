--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : c_unit.vh
--FILE GENERATED ON : Thu Aug  5 13:37:45 2010

a_unit.vhd
b_unit.vhd
c_unit.vhd
stim_expect_mem_template.vhd
tb.vhd
