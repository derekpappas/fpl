// Test type: always statement - event_trigger - no attribute instance
// Vparser rule name:
// Author: andreib
module alwcon13;
event a;
always ->a;
endmodule
