//test type : module_or_generate_item ::= module_or_generate_item_declaration (real_declaration)
//vparser rule name : 
//author : Codrin
module test_0190;
(* realnr = 1, intnr =0 *) wire out;
 assign out = 0e2;
endmodule
