// Test type: Continuous assignment - st0, wk1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous121;
wire a;
assign (strong0, weak1) a=1'b1;
endmodule
