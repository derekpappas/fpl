`include "defines.v"

module o1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 268
  output [1 - 1:0] ar_sa0_s10;
  n1 n10(.ar_sa0_s10(ar_sa0_s10));
  `include "o1.logic.vh"
endmodule

