//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : eth_mac.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module eth_mac(lbdummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 26
  input lbdummy3;
  `include "eth_mac.logic.v"
endmodule

