//test type : operator_^~ hierarchical_identifier
//vparser rule name : 
//author : Bogdan Mereghea
module unary_operator11;
    wire a, b;
    assign a = ^~b;
endmodule
