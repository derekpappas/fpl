// Test type: Decimal Numbers - upper case x digit
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'dX;
endmodule
