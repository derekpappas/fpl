// Test type: Decimal Numbers - spaces between size base and value
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=32 'd 16;
endmodule
