// Test type: Real numbers - 2 numbers
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=35.98;
endmodule
