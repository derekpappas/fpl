// Test type: Hex Numbers - no size lower case base
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a='h1A3F;
endmodule
