`ifndef DFF
`define DFF
module dff;
endmodule

module dffr;
endmodule

module dffre;
endmodule

module dffrl_async;
endmodule

module mux2ds;
endmodule

module mux3ds;
endmodule


`endif
