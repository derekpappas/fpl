/**//**/`default_nettype wire
module x;
endmodule
