// Test type: Expression - primary - hid
// Vparser rule name: 
// Author: andreib
module expressiontest;
wire a;
endmodule
