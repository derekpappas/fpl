//Primitive Instantiation and Instances: gate_instantiation = n_input_gatetype ...;
//tests by GabrielD
module gate_instantiation_n_input0;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input11;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input12;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input13;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input14;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input15;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input16;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input17;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input18;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input19;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input20;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input21;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input22;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input23;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input24;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input25;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input26;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input27;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input28;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input29;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input30;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input31;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input32;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input33;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input34;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input35;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input36;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input37;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input38;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input39;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input40;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input41;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input42;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input43;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input44;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input45;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input46;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input47;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input48;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input49;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input50;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input51;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input52;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input53;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input54;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input55;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input56;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input57;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input58;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input59;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input60;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input61;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input62;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input63;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input64;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input65;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input66;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input67;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input68;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input69;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input70;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input71;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input72;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input73;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input74;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input75;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input76;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input77;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input78;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input79;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input80;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input81;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input82;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input83;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input84;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input85;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input86;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input87;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input88;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input89;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input90;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input91;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input92;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input93;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input94;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input95;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input96;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input97;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input98;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input99;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  and (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input1999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input2999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nand (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input3999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input4999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  or (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input5999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input6999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  nor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input7999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input8999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9584;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9585;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9586;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9587;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9588;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9589;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9590;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9591;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9592;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9593;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9594;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9595;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9596;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9597;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9598;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9599;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9600;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9601;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9602;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9603;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9604;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9605;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9606;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9607;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9608;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9609;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9610;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9611;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9612;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9613;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9614;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9615;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9616;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9617;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9618;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9619;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9620;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9621;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9622;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9623;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9624;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9625;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9626;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9627;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9628;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9629;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9630;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9631;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9632;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9633;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9634;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9635;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9636;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9637;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9638;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9639;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9640;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9641;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9642;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9643;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9644;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9645;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9646;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9647;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9648;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9649;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9650;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9651;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9652;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9653;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9654;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9655;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9656;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9657;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9658;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9659;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9660;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9661;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9662;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9663;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9664;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9665;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9666;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9667;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9668;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9669;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9670;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9671;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9672;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9673;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9674;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9675;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9676;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9677;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9678;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9679;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9680;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9681;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9682;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9683;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9684;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9685;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9686;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9687;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9688;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9689;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9690;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9691;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9692;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9693;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9694;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9695;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9696;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9697;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9698;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9699;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9700;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9701;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9702;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9703;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9704;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9705;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9706;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9707;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9708;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9709;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9710;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9711;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9712;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9713;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9714;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9715;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9716;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9717;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9718;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9719;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9720;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9721;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9722;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9723;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9724;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9725;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9726;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9727;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9728;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9729;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9730;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9731;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9732;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9733;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9734;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9735;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9736;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9737;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9738;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9739;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9740;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9741;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9742;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9743;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9744;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9745;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9746;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9747;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9748;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9749;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9750;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9751;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9752;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9753;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9754;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9755;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9756;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9757;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9758;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9759;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9760;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9761;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9762;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9763;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9764;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9765;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9766;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9767;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9768;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9769;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9770;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9771;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9772;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9773;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9774;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9775;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9776;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9777;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9778;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9779;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9780;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9781;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9782;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9783;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9784;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9785;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9786;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9787;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9788;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9789;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9790;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9791;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9792;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9793;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9794;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9795;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9796;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9797;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9798;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9799;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9800;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9801;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9802;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9803;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9804;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9805;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9806;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9807;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9808;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9809;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9810;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9811;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9812;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9813;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9814;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9815;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9816;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9817;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9818;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9819;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9820;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9821;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9822;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9823;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9824;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9825;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9826;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9827;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9828;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9829;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9830;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9831;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9832;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9833;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9834;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9835;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9836;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9837;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9838;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9839;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9840;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9841;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9842;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9843;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9844;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9845;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9846;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9847;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9848;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9849;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9850;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9851;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9852;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9853;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9854;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9855;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9856;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9857;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9858;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9859;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9860;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9861;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9862;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9863;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9864;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9865;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9866;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9867;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9868;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9869;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9870;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9871;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9872;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9873;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9874;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9875;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9876;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9877;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9878;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9879;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9880;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9881;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9882;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9883;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9884;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9885;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9886;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9887;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9888;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9889;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9890;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9891;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9892;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9893;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9894;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9895;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9896;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9897;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9898;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9899;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9900;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9901;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9902;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9903;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9904;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9905;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9906;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9907;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9908;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9909;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9910;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9911;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9912;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9913;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9914;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9915;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9916;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9917;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9918;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9919;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9920;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9921;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9922;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9923;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9924;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9925;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9926;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9927;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9928;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9929;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9930;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9931;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9932;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9933;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9934;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9935;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9936;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9937;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9938;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9939;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9940;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9941;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9942;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9943;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9944;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9945;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9946;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9947;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9948;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9949;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9950;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9951;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9952;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9953;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9954;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9955;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9956;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9957;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9958;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9959;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9960;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9961;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9962;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9963;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9964;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9965;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9966;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9967;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9968;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9969;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9970;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9971;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9972;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9973;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9974;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9975;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9976;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9977;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9978;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9979;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9980;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9981;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9982;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9983;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9984;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9985;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9986;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9987;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9988;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9989;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9990;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9991;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9992;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9993;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9994;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9995;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (highz0,strong1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9996;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9997;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9998;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input9999;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10000;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10001;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10002;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10003;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10004;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10005;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10006;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10007;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10008;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10009;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10010;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10011;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10012;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10013;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10014;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10015;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10016;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10017;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10018;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10019;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10020;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10021;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10022;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10023;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10024;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10025;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10026;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10027;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10028;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10029;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10030;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10031;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10032;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10033;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10034;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10035;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10036;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10037;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10038;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10039;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10040;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10041;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10042;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10043;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10044;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10045;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10046;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10047;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10048;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10049;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10050;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10051;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10052;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10053;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10054;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10055;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10056;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10057;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10058;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10059;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10060;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10061;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10062;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10063;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10064;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10065;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10066;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10067;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10068;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10069;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10070;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10071;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10072;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10073;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10074;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10075;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10076;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10077;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10078;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10079;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10080;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10081;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10082;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10083;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10084;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10085;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10086;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10087;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10088;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10089;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10090;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10091;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10092;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10093;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10094;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10095;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10096;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10097;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10098;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10099;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10100;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10101;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10102;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10103;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10104;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10105;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10106;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10107;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10108;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10109;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10110;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10111;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10112;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10113;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10114;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10115;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10116;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10117;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10118;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10119;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10120;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10121;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10122;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10123;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10124;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10125;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10126;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10127;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10128;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10129;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10130;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10131;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10132;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10133;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10134;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10135;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10136;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10137;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10138;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10139;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10140;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10141;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10142;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10143;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10144;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10145;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10146;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10147;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10148;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10149;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10150;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10151;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10152;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10153;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10154;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10155;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10156;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10157;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10158;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10159;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10160;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10161;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10162;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10163;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10164;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10165;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10166;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10167;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10168;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10169;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10170;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10171;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10172;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10173;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10174;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10175;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10176;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10177;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10178;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10179;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10180;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10181;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10182;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10183;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10184;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10185;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10186;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10187;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10188;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10189;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10190;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10191;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10192;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10193;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10194;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10195;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10196;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10197;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10198;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10199;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10200;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10201;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10202;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10203;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10204;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10205;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10206;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10207;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10208;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10209;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10210;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10211;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10212;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10213;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10214;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10215;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10216;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10217;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10218;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10219;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10220;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10221;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10222;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10223;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10224;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10225;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10226;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10227;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10228;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10229;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10230;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10231;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10232;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10233;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10234;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10235;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10236;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10237;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10238;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10239;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10240;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10241;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10242;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10243;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10244;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10245;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10246;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10247;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10248;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10249;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10250;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10251;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10252;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10253;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10254;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10255;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10256;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10257;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10258;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10259;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10260;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10261;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10262;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10263;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10264;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10265;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10266;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10267;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10268;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10269;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10270;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10271;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10272;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10273;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10274;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10275;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10276;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10277;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10278;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10279;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10280;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10281;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10282;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10283;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10284;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10285;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10286;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10287;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10288;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10289;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10290;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10291;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10292;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10293;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10294;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10295;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10296;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10297;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10298;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10299;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10300;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10301;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10302;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10303;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10304;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10305;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10306;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10307;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10308;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10309;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10310;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10311;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10312;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10313;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10314;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10315;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10316;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10317;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10318;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10319;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10320;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10321;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10322;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10323;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10324;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10325;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10326;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10327;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10328;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10329;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10330;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10331;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10332;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10333;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10334;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10335;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10336;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10337;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10338;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10339;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10340;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10341;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10342;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10343;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10344;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10345;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10346;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10347;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10348;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10349;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10350;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10351;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10352;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10353;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10354;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10355;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10356;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10357;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10358;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10359;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10360;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10361;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10362;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10363;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10364;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10365;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10366;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10367;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10368;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10369;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10370;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10371;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10372;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10373;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10374;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10375;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10376;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10377;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10378;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10379;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10380;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10381;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10382;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10383;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10384;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10385;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10386;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10387;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10388;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10389;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10390;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10391;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10392;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10393;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10394;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10395;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10396;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10397;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10398;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10399;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10400;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10401;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10402;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10403;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10404;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10405;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10406;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10407;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10408;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10409;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10410;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10411;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10412;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10413;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10414;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10415;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10416;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10417;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10418;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10419;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10420;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10421;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10422;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10423;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10424;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10425;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10426;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10427;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10428;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10429;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10430;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10431;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10432;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10433;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10434;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10435;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10436;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10437;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10438;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10439;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10440;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10441;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10442;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10443;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10444;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10445;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10446;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10447;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10448;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10449;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10450;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10451;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10452;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10453;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10454;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10455;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10456;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10457;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10458;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10459;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10460;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10461;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10462;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10463;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10464;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10465;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10466;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10467;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10468;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10469;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10470;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10471;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10472;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10473;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10474;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10475;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10476;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10477;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10478;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10479;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10480;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10481;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10482;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10483;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10484;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10485;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10486;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10487;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10488;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10489;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10490;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10491;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10492;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10493;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10494;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10495;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10496;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10497;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10498;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10499;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10500;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10501;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10502;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10503;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10504;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10505;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10506;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10507;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10508;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10509;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10510;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10511;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10512;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10513;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10514;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10515;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10516;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10517;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10518;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10519;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10520;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10521;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10522;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10523;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10524;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10525;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10526;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10527;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10528;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10529;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10530;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10531;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10532;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10533;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10534;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10535;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10536;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10537;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10538;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10539;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10540;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10541;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10542;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10543;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10544;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10545;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10546;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10547;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10548;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10549;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10550;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10551;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10552;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10553;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10554;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10555;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10556;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10557;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10558;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10559;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10560;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10561;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10562;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10563;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10564;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10565;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10566;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10567;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10568;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10569;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10570;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10571;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10572;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10573;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10574;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10575;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10576;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10577;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10578;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10579;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10580;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10581;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10582;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ) ;
endmodule
module gate_instantiation_n_input10583;
  wire output_terminal, ncontrol_terminal;
  reg input_terminal, pcontrol_terminal;
  xnor (supply0,highz1) #2 name1 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name2 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) , name3 (output_terminal ,input_terminal ,input_terminal ,input_terminal ,input_terminal ) ;
endmodule
