module x;

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify
specify endspecify

endmodule
