// Test type: initial statement - system_task_enable - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon34;
reg a;
initial a=$random;
endmodule
