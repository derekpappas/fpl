//test type : port_declaration
//vparser rule name : 
//author : Codrin
module declaration_0140(x);
 (* a = 5, b = 11 *) inout x;
endmodule
