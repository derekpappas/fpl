// Test type: Continuous assignment - h0, sup1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous616;
wire a;
assign (highz0, supply1) a=1'b1;
endmodule
