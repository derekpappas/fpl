`include "defines.v"

module crcr();
// Location of source csl unit: file name = IPX2400.csl line number = 56
  `include "crcr.logic.v"
endmodule

