module testbench_input_declaration;
    input_declaration0 input_declaration_instance0();
    input_declaration1 input_declaration_instance1();
    input_declaration2 input_declaration_instance2();
    input_declaration3 input_declaration_instance3();
    input_declaration4 input_declaration_instance4();
    input_declaration5 input_declaration_instance5();
    input_declaration6 input_declaration_instance6();
    input_declaration7 input_declaration_instance7();
    input_declaration8 input_declaration_instance8();
    input_declaration9 input_declaration_instance9();
    input_declaration10 input_declaration_instance10();
    input_declaration11 input_declaration_instance11();
    input_declaration12 input_declaration_instance12();
    input_declaration13 input_declaration_instance13();
    input_declaration14 input_declaration_instance14();
    input_declaration15 input_declaration_instance15();
    input_declaration16 input_declaration_instance16();
    input_declaration17 input_declaration_instance17();
    input_declaration18 input_declaration_instance18();
    input_declaration19 input_declaration_instance19();
    input_declaration20 input_declaration_instance20();
    input_declaration21 input_declaration_instance21();
    input_declaration22 input_declaration_instance22();
    input_declaration23 input_declaration_instance23();
    input_declaration24 input_declaration_instance24();
    input_declaration25 input_declaration_instance25();
    input_declaration26 input_declaration_instance26();
    input_declaration27 input_declaration_instance27();
    input_declaration28 input_declaration_instance28();
    input_declaration29 input_declaration_instance29();
    input_declaration30 input_declaration_instance30();
    input_declaration31 input_declaration_instance31();
    input_declaration32 input_declaration_instance32();
    input_declaration33 input_declaration_instance33();
    input_declaration34 input_declaration_instance34();
    input_declaration35 input_declaration_instance35();
    input_declaration36 input_declaration_instance36();
    input_declaration37 input_declaration_instance37();
    input_declaration38 input_declaration_instance38();
    input_declaration39 input_declaration_instance39();
    input_declaration40 input_declaration_instance40();
    input_declaration41 input_declaration_instance41();
    input_declaration42 input_declaration_instance42();
    input_declaration43 input_declaration_instance43();
    input_declaration44 input_declaration_instance44();
    input_declaration45 input_declaration_instance45();
    input_declaration46 input_declaration_instance46();
    input_declaration47 input_declaration_instance47();
    input_declaration48 input_declaration_instance48();
    input_declaration49 input_declaration_instance49();
    input_declaration50 input_declaration_instance50();
    input_declaration51 input_declaration_instance51();
    input_declaration52 input_declaration_instance52();
    input_declaration53 input_declaration_instance53();
    input_declaration54 input_declaration_instance54();
    input_declaration55 input_declaration_instance55();
    input_declaration56 input_declaration_instance56();
    input_declaration57 input_declaration_instance57();
    input_declaration58 input_declaration_instance58();
    input_declaration59 input_declaration_instance59();
    input_declaration60 input_declaration_instance60();
    input_declaration61 input_declaration_instance61();
    input_declaration62 input_declaration_instance62();
    input_declaration63 input_declaration_instance63();
    input_declaration64 input_declaration_instance64();
    input_declaration65 input_declaration_instance65();
    input_declaration66 input_declaration_instance66();
    input_declaration67 input_declaration_instance67();
    input_declaration68 input_declaration_instance68();
    input_declaration69 input_declaration_instance69();
    input_declaration70 input_declaration_instance70();
    input_declaration71 input_declaration_instance71();
    input_declaration72 input_declaration_instance72();
    input_declaration73 input_declaration_instance73();
    input_declaration74 input_declaration_instance74();
    input_declaration75 input_declaration_instance75();
    input_declaration76 input_declaration_instance76();
    input_declaration77 input_declaration_instance77();
    input_declaration78 input_declaration_instance78();
    input_declaration79 input_declaration_instance79();
    input_declaration80 input_declaration_instance80();
    input_declaration81 input_declaration_instance81();
    input_declaration82 input_declaration_instance82();
    input_declaration83 input_declaration_instance83();
    input_declaration84 input_declaration_instance84();
    input_declaration85 input_declaration_instance85();
    input_declaration86 input_declaration_instance86();
    input_declaration87 input_declaration_instance87();
    input_declaration88 input_declaration_instance88();
    input_declaration89 input_declaration_instance89();
    input_declaration90 input_declaration_instance90();
    input_declaration91 input_declaration_instance91();
    input_declaration92 input_declaration_instance92();
    input_declaration93 input_declaration_instance93();
    input_declaration94 input_declaration_instance94();
    input_declaration95 input_declaration_instance95();
    input_declaration96 input_declaration_instance96();
    input_declaration97 input_declaration_instance97();
    input_declaration98 input_declaration_instance98();
    input_declaration99 input_declaration_instance99();
    input_declaration100 input_declaration_instance100();
    input_declaration101 input_declaration_instance101();
    input_declaration102 input_declaration_instance102();
    input_declaration103 input_declaration_instance103();
    input_declaration104 input_declaration_instance104();
    input_declaration105 input_declaration_instance105();
    input_declaration106 input_declaration_instance106();
    input_declaration107 input_declaration_instance107();
    input_declaration108 input_declaration_instance108();
    input_declaration109 input_declaration_instance109();
    input_declaration110 input_declaration_instance110();
    input_declaration111 input_declaration_instance111();
    input_declaration112 input_declaration_instance112();
    input_declaration113 input_declaration_instance113();
    input_declaration114 input_declaration_instance114();
    input_declaration115 input_declaration_instance115();
    input_declaration116 input_declaration_instance116();
    input_declaration117 input_declaration_instance117();
    input_declaration118 input_declaration_instance118();
    input_declaration119 input_declaration_instance119();
    input_declaration120 input_declaration_instance120();
    input_declaration121 input_declaration_instance121();
    input_declaration122 input_declaration_instance122();
    input_declaration123 input_declaration_instance123();
    input_declaration124 input_declaration_instance124();
    input_declaration125 input_declaration_instance125();
    input_declaration126 input_declaration_instance126();
    input_declaration127 input_declaration_instance127();
    input_declaration128 input_declaration_instance128();
    input_declaration129 input_declaration_instance129();
    input_declaration130 input_declaration_instance130();
    input_declaration131 input_declaration_instance131();
    input_declaration132 input_declaration_instance132();
    input_declaration133 input_declaration_instance133();
    input_declaration134 input_declaration_instance134();
    input_declaration135 input_declaration_instance135();
    input_declaration136 input_declaration_instance136();
    input_declaration137 input_declaration_instance137();
    input_declaration138 input_declaration_instance138();
    input_declaration139 input_declaration_instance139();
    input_declaration140 input_declaration_instance140();
    input_declaration141 input_declaration_instance141();
    input_declaration142 input_declaration_instance142();
    input_declaration143 input_declaration_instance143();
    input_declaration144 input_declaration_instance144();
    input_declaration145 input_declaration_instance145();
    input_declaration146 input_declaration_instance146();
    input_declaration147 input_declaration_instance147();
    input_declaration148 input_declaration_instance148();
    input_declaration149 input_declaration_instance149();
    input_declaration150 input_declaration_instance150();
    input_declaration151 input_declaration_instance151();
    input_declaration152 input_declaration_instance152();
    input_declaration153 input_declaration_instance153();
    input_declaration154 input_declaration_instance154();
    input_declaration155 input_declaration_instance155();
    input_declaration156 input_declaration_instance156();
    input_declaration157 input_declaration_instance157();
    input_declaration158 input_declaration_instance158();
    input_declaration159 input_declaration_instance159();
    input_declaration160 input_declaration_instance160();
    input_declaration161 input_declaration_instance161();
    input_declaration162 input_declaration_instance162();
    input_declaration163 input_declaration_instance163();
    input_declaration164 input_declaration_instance164();
    input_declaration165 input_declaration_instance165();
    input_declaration166 input_declaration_instance166();
    input_declaration167 input_declaration_instance167();
    input_declaration168 input_declaration_instance168();
    input_declaration169 input_declaration_instance169();
    input_declaration170 input_declaration_instance170();
    input_declaration171 input_declaration_instance171();
    input_declaration172 input_declaration_instance172();
    input_declaration173 input_declaration_instance173();
    input_declaration174 input_declaration_instance174();
    input_declaration175 input_declaration_instance175();
    input_declaration176 input_declaration_instance176();
    input_declaration177 input_declaration_instance177();
    input_declaration178 input_declaration_instance178();
    input_declaration179 input_declaration_instance179();
    input_declaration180 input_declaration_instance180();
    input_declaration181 input_declaration_instance181();
    input_declaration182 input_declaration_instance182();
    input_declaration183 input_declaration_instance183();
    input_declaration184 input_declaration_instance184();
    input_declaration185 input_declaration_instance185();
    input_declaration186 input_declaration_instance186();
    input_declaration187 input_declaration_instance187();
    input_declaration188 input_declaration_instance188();
    input_declaration189 input_declaration_instance189();
    input_declaration190 input_declaration_instance190();
    input_declaration191 input_declaration_instance191();
    input_declaration192 input_declaration_instance192();
    input_declaration193 input_declaration_instance193();
    input_declaration194 input_declaration_instance194();
    input_declaration195 input_declaration_instance195();
    input_declaration196 input_declaration_instance196();
    input_declaration197 input_declaration_instance197();
    input_declaration198 input_declaration_instance198();
    input_declaration199 input_declaration_instance199();
    input_declaration200 input_declaration_instance200();
    input_declaration201 input_declaration_instance201();
    input_declaration202 input_declaration_instance202();
    input_declaration203 input_declaration_instance203();
    input_declaration204 input_declaration_instance204();
    input_declaration205 input_declaration_instance205();
    input_declaration206 input_declaration_instance206();
    input_declaration207 input_declaration_instance207();
    input_declaration208 input_declaration_instance208();
    input_declaration209 input_declaration_instance209();
    input_declaration210 input_declaration_instance210();
    input_declaration211 input_declaration_instance211();
    input_declaration212 input_declaration_instance212();
    input_declaration213 input_declaration_instance213();
    input_declaration214 input_declaration_instance214();
    input_declaration215 input_declaration_instance215();
    input_declaration216 input_declaration_instance216();
    input_declaration217 input_declaration_instance217();
    input_declaration218 input_declaration_instance218();
    input_declaration219 input_declaration_instance219();
    input_declaration220 input_declaration_instance220();
    input_declaration221 input_declaration_instance221();
    input_declaration222 input_declaration_instance222();
    input_declaration223 input_declaration_instance223();
    input_declaration224 input_declaration_instance224();
    input_declaration225 input_declaration_instance225();
    input_declaration226 input_declaration_instance226();
    input_declaration227 input_declaration_instance227();
    input_declaration228 input_declaration_instance228();
    input_declaration229 input_declaration_instance229();
    input_declaration230 input_declaration_instance230();
    input_declaration231 input_declaration_instance231();
    input_declaration232 input_declaration_instance232();
    input_declaration233 input_declaration_instance233();
    input_declaration234 input_declaration_instance234();
    input_declaration235 input_declaration_instance235();
    input_declaration236 input_declaration_instance236();
    input_declaration237 input_declaration_instance237();
    input_declaration238 input_declaration_instance238();
    input_declaration239 input_declaration_instance239();
    input_declaration240 input_declaration_instance240();
    input_declaration241 input_declaration_instance241();
    input_declaration242 input_declaration_instance242();
    input_declaration243 input_declaration_instance243();
    input_declaration244 input_declaration_instance244();
    input_declaration245 input_declaration_instance245();
    input_declaration246 input_declaration_instance246();
    input_declaration247 input_declaration_instance247();
    input_declaration248 input_declaration_instance248();
    input_declaration249 input_declaration_instance249();
    input_declaration250 input_declaration_instance250();
    input_declaration251 input_declaration_instance251();
    input_declaration252 input_declaration_instance252();
    input_declaration253 input_declaration_instance253();
    input_declaration254 input_declaration_instance254();
    input_declaration255 input_declaration_instance255();
    input_declaration256 input_declaration_instance256();
    input_declaration257 input_declaration_instance257();
    input_declaration258 input_declaration_instance258();
    input_declaration259 input_declaration_instance259();
    input_declaration260 input_declaration_instance260();
    input_declaration261 input_declaration_instance261();
    input_declaration262 input_declaration_instance262();
    input_declaration263 input_declaration_instance263();
    input_declaration264 input_declaration_instance264();
    input_declaration265 input_declaration_instance265();
    input_declaration266 input_declaration_instance266();
    input_declaration267 input_declaration_instance267();
    input_declaration268 input_declaration_instance268();
    input_declaration269 input_declaration_instance269();
    input_declaration270 input_declaration_instance270();
    input_declaration271 input_declaration_instance271();
    input_declaration272 input_declaration_instance272();
    input_declaration273 input_declaration_instance273();
    input_declaration274 input_declaration_instance274();
    input_declaration275 input_declaration_instance275();
    input_declaration276 input_declaration_instance276();
    input_declaration277 input_declaration_instance277();
    input_declaration278 input_declaration_instance278();
    input_declaration279 input_declaration_instance279();
    input_declaration280 input_declaration_instance280();
    input_declaration281 input_declaration_instance281();
    input_declaration282 input_declaration_instance282();
    input_declaration283 input_declaration_instance283();
    input_declaration284 input_declaration_instance284();
    input_declaration285 input_declaration_instance285();
    input_declaration286 input_declaration_instance286();
    input_declaration287 input_declaration_instance287();
    input_declaration288 input_declaration_instance288();
    input_declaration289 input_declaration_instance289();
    input_declaration290 input_declaration_instance290();
    input_declaration291 input_declaration_instance291();
    input_declaration292 input_declaration_instance292();
    input_declaration293 input_declaration_instance293();
    input_declaration294 input_declaration_instance294();
    input_declaration295 input_declaration_instance295();
    input_declaration296 input_declaration_instance296();
    input_declaration297 input_declaration_instance297();
    input_declaration298 input_declaration_instance298();
    input_declaration299 input_declaration_instance299();
    input_declaration300 input_declaration_instance300();
    input_declaration301 input_declaration_instance301();
    input_declaration302 input_declaration_instance302();
    input_declaration303 input_declaration_instance303();
    input_declaration304 input_declaration_instance304();
    input_declaration305 input_declaration_instance305();
    input_declaration306 input_declaration_instance306();
    input_declaration307 input_declaration_instance307();
    input_declaration308 input_declaration_instance308();
    input_declaration309 input_declaration_instance309();
    input_declaration310 input_declaration_instance310();
    input_declaration311 input_declaration_instance311();
    input_declaration312 input_declaration_instance312();
    input_declaration313 input_declaration_instance313();
    input_declaration314 input_declaration_instance314();
    input_declaration315 input_declaration_instance315();
    input_declaration316 input_declaration_instance316();
    input_declaration317 input_declaration_instance317();
    input_declaration318 input_declaration_instance318();
    input_declaration319 input_declaration_instance319();
    input_declaration320 input_declaration_instance320();
    input_declaration321 input_declaration_instance321();
    input_declaration322 input_declaration_instance322();
    input_declaration323 input_declaration_instance323();
    input_declaration324 input_declaration_instance324();
    input_declaration325 input_declaration_instance325();
    input_declaration326 input_declaration_instance326();
    input_declaration327 input_declaration_instance327();
    input_declaration328 input_declaration_instance328();
    input_declaration329 input_declaration_instance329();
    input_declaration330 input_declaration_instance330();
    input_declaration331 input_declaration_instance331();
    input_declaration332 input_declaration_instance332();
    input_declaration333 input_declaration_instance333();
    input_declaration334 input_declaration_instance334();
    input_declaration335 input_declaration_instance335();
    input_declaration336 input_declaration_instance336();
    input_declaration337 input_declaration_instance337();
    input_declaration338 input_declaration_instance338();
    input_declaration339 input_declaration_instance339();
    input_declaration340 input_declaration_instance340();
    input_declaration341 input_declaration_instance341();
    input_declaration342 input_declaration_instance342();
    input_declaration343 input_declaration_instance343();
    input_declaration344 input_declaration_instance344();
    input_declaration345 input_declaration_instance345();
    input_declaration346 input_declaration_instance346();
    input_declaration347 input_declaration_instance347();
    input_declaration348 input_declaration_instance348();
    input_declaration349 input_declaration_instance349();
    input_declaration350 input_declaration_instance350();
    input_declaration351 input_declaration_instance351();
    input_declaration352 input_declaration_instance352();
    input_declaration353 input_declaration_instance353();
    input_declaration354 input_declaration_instance354();
    input_declaration355 input_declaration_instance355();
    input_declaration356 input_declaration_instance356();
    input_declaration357 input_declaration_instance357();
    input_declaration358 input_declaration_instance358();
    input_declaration359 input_declaration_instance359();
    input_declaration360 input_declaration_instance360();
    input_declaration361 input_declaration_instance361();
    input_declaration362 input_declaration_instance362();
    input_declaration363 input_declaration_instance363();
    input_declaration364 input_declaration_instance364();
    input_declaration365 input_declaration_instance365();
    input_declaration366 input_declaration_instance366();
    input_declaration367 input_declaration_instance367();
    input_declaration368 input_declaration_instance368();
    input_declaration369 input_declaration_instance369();
    input_declaration370 input_declaration_instance370();
    input_declaration371 input_declaration_instance371();
    input_declaration372 input_declaration_instance372();
    input_declaration373 input_declaration_instance373();
    input_declaration374 input_declaration_instance374();
    input_declaration375 input_declaration_instance375();
    input_declaration376 input_declaration_instance376();
    input_declaration377 input_declaration_instance377();
    input_declaration378 input_declaration_instance378();
    input_declaration379 input_declaration_instance379();
    input_declaration380 input_declaration_instance380();
    input_declaration381 input_declaration_instance381();
    input_declaration382 input_declaration_instance382();
    input_declaration383 input_declaration_instance383();
    input_declaration384 input_declaration_instance384();
    input_declaration385 input_declaration_instance385();
    input_declaration386 input_declaration_instance386();
    input_declaration387 input_declaration_instance387();
    input_declaration388 input_declaration_instance388();
    input_declaration389 input_declaration_instance389();
    input_declaration390 input_declaration_instance390();
    input_declaration391 input_declaration_instance391();
    input_declaration392 input_declaration_instance392();
    input_declaration393 input_declaration_instance393();
    input_declaration394 input_declaration_instance394();
    input_declaration395 input_declaration_instance395();
    input_declaration396 input_declaration_instance396();
    input_declaration397 input_declaration_instance397();
    input_declaration398 input_declaration_instance398();
    input_declaration399 input_declaration_instance399();
    input_declaration400 input_declaration_instance400();
    input_declaration401 input_declaration_instance401();
    input_declaration402 input_declaration_instance402();
    input_declaration403 input_declaration_instance403();
    input_declaration404 input_declaration_instance404();
    input_declaration405 input_declaration_instance405();
    input_declaration406 input_declaration_instance406();
    input_declaration407 input_declaration_instance407();
    input_declaration408 input_declaration_instance408();
    input_declaration409 input_declaration_instance409();
    input_declaration410 input_declaration_instance410();
    input_declaration411 input_declaration_instance411();
    input_declaration412 input_declaration_instance412();
    input_declaration413 input_declaration_instance413();
    input_declaration414 input_declaration_instance414();
    input_declaration415 input_declaration_instance415();
    input_declaration416 input_declaration_instance416();
    input_declaration417 input_declaration_instance417();
    input_declaration418 input_declaration_instance418();
    input_declaration419 input_declaration_instance419();
    input_declaration420 input_declaration_instance420();
    input_declaration421 input_declaration_instance421();
    input_declaration422 input_declaration_instance422();
    input_declaration423 input_declaration_instance423();
    input_declaration424 input_declaration_instance424();
    input_declaration425 input_declaration_instance425();
    input_declaration426 input_declaration_instance426();
    input_declaration427 input_declaration_instance427();
    input_declaration428 input_declaration_instance428();
    input_declaration429 input_declaration_instance429();
    input_declaration430 input_declaration_instance430();
    input_declaration431 input_declaration_instance431();
    input_declaration432 input_declaration_instance432();
    input_declaration433 input_declaration_instance433();
    input_declaration434 input_declaration_instance434();
    input_declaration435 input_declaration_instance435();
    input_declaration436 input_declaration_instance436();
    input_declaration437 input_declaration_instance437();
    input_declaration438 input_declaration_instance438();
    input_declaration439 input_declaration_instance439();
    input_declaration440 input_declaration_instance440();
    input_declaration441 input_declaration_instance441();
    input_declaration442 input_declaration_instance442();
    input_declaration443 input_declaration_instance443();
    input_declaration444 input_declaration_instance444();
    input_declaration445 input_declaration_instance445();
    input_declaration446 input_declaration_instance446();
    input_declaration447 input_declaration_instance447();
    input_declaration448 input_declaration_instance448();
    input_declaration449 input_declaration_instance449();
    input_declaration450 input_declaration_instance450();
    input_declaration451 input_declaration_instance451();
    input_declaration452 input_declaration_instance452();
    input_declaration453 input_declaration_instance453();
    input_declaration454 input_declaration_instance454();
    input_declaration455 input_declaration_instance455();
    input_declaration456 input_declaration_instance456();
    input_declaration457 input_declaration_instance457();
    input_declaration458 input_declaration_instance458();
    input_declaration459 input_declaration_instance459();
    input_declaration460 input_declaration_instance460();
    input_declaration461 input_declaration_instance461();
    input_declaration462 input_declaration_instance462();
    input_declaration463 input_declaration_instance463();
    input_declaration464 input_declaration_instance464();
    input_declaration465 input_declaration_instance465();
    input_declaration466 input_declaration_instance466();
    input_declaration467 input_declaration_instance467();
    input_declaration468 input_declaration_instance468();
    input_declaration469 input_declaration_instance469();
    input_declaration470 input_declaration_instance470();
    input_declaration471 input_declaration_instance471();
    input_declaration472 input_declaration_instance472();
    input_declaration473 input_declaration_instance473();
    input_declaration474 input_declaration_instance474();
    input_declaration475 input_declaration_instance475();
    input_declaration476 input_declaration_instance476();
    input_declaration477 input_declaration_instance477();
    input_declaration478 input_declaration_instance478();
    input_declaration479 input_declaration_instance479();
    input_declaration480 input_declaration_instance480();
    input_declaration481 input_declaration_instance481();
    input_declaration482 input_declaration_instance482();
    input_declaration483 input_declaration_instance483();
    input_declaration484 input_declaration_instance484();
    input_declaration485 input_declaration_instance485();
    input_declaration486 input_declaration_instance486();
    input_declaration487 input_declaration_instance487();
    input_declaration488 input_declaration_instance488();
    input_declaration489 input_declaration_instance489();
    input_declaration490 input_declaration_instance490();
    input_declaration491 input_declaration_instance491();
    input_declaration492 input_declaration_instance492();
    input_declaration493 input_declaration_instance493();
    input_declaration494 input_declaration_instance494();
    input_declaration495 input_declaration_instance495();
    input_declaration496 input_declaration_instance496();
    input_declaration497 input_declaration_instance497();
    input_declaration498 input_declaration_instance498();
    input_declaration499 input_declaration_instance499();
    input_declaration500 input_declaration_instance500();
    input_declaration501 input_declaration_instance501();
    input_declaration502 input_declaration_instance502();
    input_declaration503 input_declaration_instance503();
    input_declaration504 input_declaration_instance504();
    input_declaration505 input_declaration_instance505();
    input_declaration506 input_declaration_instance506();
    input_declaration507 input_declaration_instance507();
    input_declaration508 input_declaration_instance508();
    input_declaration509 input_declaration_instance509();
    input_declaration510 input_declaration_instance510();
    input_declaration511 input_declaration_instance511();
    input_declaration512 input_declaration_instance512();
    input_declaration513 input_declaration_instance513();
    input_declaration514 input_declaration_instance514();
    input_declaration515 input_declaration_instance515();
    input_declaration516 input_declaration_instance516();
    input_declaration517 input_declaration_instance517();
    input_declaration518 input_declaration_instance518();
    input_declaration519 input_declaration_instance519();
    input_declaration520 input_declaration_instance520();
    input_declaration521 input_declaration_instance521();
    input_declaration522 input_declaration_instance522();
    input_declaration523 input_declaration_instance523();
    input_declaration524 input_declaration_instance524();
    input_declaration525 input_declaration_instance525();
    input_declaration526 input_declaration_instance526();
    input_declaration527 input_declaration_instance527();
    input_declaration528 input_declaration_instance528();
    input_declaration529 input_declaration_instance529();
    input_declaration530 input_declaration_instance530();
    input_declaration531 input_declaration_instance531();
    input_declaration532 input_declaration_instance532();
    input_declaration533 input_declaration_instance533();
    input_declaration534 input_declaration_instance534();
    input_declaration535 input_declaration_instance535();
    input_declaration536 input_declaration_instance536();
    input_declaration537 input_declaration_instance537();
    input_declaration538 input_declaration_instance538();
    input_declaration539 input_declaration_instance539();
    input_declaration540 input_declaration_instance540();
    input_declaration541 input_declaration_instance541();
    input_declaration542 input_declaration_instance542();
    input_declaration543 input_declaration_instance543();
    input_declaration544 input_declaration_instance544();
    input_declaration545 input_declaration_instance545();
    input_declaration546 input_declaration_instance546();
    input_declaration547 input_declaration_instance547();
    input_declaration548 input_declaration_instance548();
    input_declaration549 input_declaration_instance549();
    input_declaration550 input_declaration_instance550();
    input_declaration551 input_declaration_instance551();
    input_declaration552 input_declaration_instance552();
    input_declaration553 input_declaration_instance553();
    input_declaration554 input_declaration_instance554();
    input_declaration555 input_declaration_instance555();
    input_declaration556 input_declaration_instance556();
    input_declaration557 input_declaration_instance557();
    input_declaration558 input_declaration_instance558();
    input_declaration559 input_declaration_instance559();
    input_declaration560 input_declaration_instance560();
    input_declaration561 input_declaration_instance561();
    input_declaration562 input_declaration_instance562();
    input_declaration563 input_declaration_instance563();
    input_declaration564 input_declaration_instance564();
    input_declaration565 input_declaration_instance565();
    input_declaration566 input_declaration_instance566();
    input_declaration567 input_declaration_instance567();
    input_declaration568 input_declaration_instance568();
    input_declaration569 input_declaration_instance569();
    input_declaration570 input_declaration_instance570();
    input_declaration571 input_declaration_instance571();
endmodule
//@
//author : andreib
module input_declaration0( abc,ABC ); input abc,ABC;
endmodule
//author : andreib
module input_declaration1( abc,ABC ); input [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration2( abc,ABC ); input [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration3( abc,ABC ); input [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration4( abc,ABC ); input [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration5( abc,ABC ); input [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration6( abc,ABC ); input [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration7( abc,ABC ); input [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration8( abc,ABC ); input [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration9( abc,ABC ); input [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration10( abc,ABC ); input [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration11( abc,ABC ); input [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration12( abc,ABC ); input [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration13( abc,ABC ); input [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration14( abc,ABC ); input [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration15( abc,ABC ); input [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration16( abc,ABC ); input [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration17( abc,ABC ); input [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration18( abc,ABC ); input [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration19( abc,ABC ); input [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration20( abc,ABC ); input [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration21( abc,ABC ); input [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration22( abc,ABC ); input [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration23( abc,ABC ); input [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration24( abc,ABC ); input [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration25( abc,ABC ); input [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration26( abc,ABC ); input signed abc,ABC;
endmodule
//author : andreib
module input_declaration27( abc,ABC ); input signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration28( abc,ABC ); input signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration29( abc,ABC ); input signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration30( abc,ABC ); input signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration31( abc,ABC ); input signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration32( abc,ABC ); input signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration33( abc,ABC ); input signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration34( abc,ABC ); input signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration35( abc,ABC ); input signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration36( abc,ABC ); input signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration37( abc,ABC ); input signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration38( abc,ABC ); input signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration39( abc,ABC ); input signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration40( abc,ABC ); input signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration41( abc,ABC ); input signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration42( abc,ABC ); input signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration43( abc,ABC ); input signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration44( abc,ABC ); input signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration45( abc,ABC ); input signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration46( abc,ABC ); input signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration47( abc,ABC ); input signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration48( abc,ABC ); input signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration49( abc,ABC ); input signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration50( abc,ABC ); input signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration51( abc,ABC ); input signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration52( abc,ABC ); input supply0 abc,ABC;
endmodule
//author : andreib
module input_declaration53( abc,ABC ); input supply0 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration54( abc,ABC ); input supply0 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration55( abc,ABC ); input supply0 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration56( abc,ABC ); input supply0 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration57( abc,ABC ); input supply0 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration58( abc,ABC ); input supply0 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration59( abc,ABC ); input supply0 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration60( abc,ABC ); input supply0 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration61( abc,ABC ); input supply0 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration62( abc,ABC ); input supply0 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration63( abc,ABC ); input supply0 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration64( abc,ABC ); input supply0 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration65( abc,ABC ); input supply0 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration66( abc,ABC ); input supply0 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration67( abc,ABC ); input supply0 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration68( abc,ABC ); input supply0 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration69( abc,ABC ); input supply0 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration70( abc,ABC ); input supply0 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration71( abc,ABC ); input supply0 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration72( abc,ABC ); input supply0 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration73( abc,ABC ); input supply0 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration74( abc,ABC ); input supply0 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration75( abc,ABC ); input supply0 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration76( abc,ABC ); input supply0 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration77( abc,ABC ); input supply0 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration78( abc,ABC ); input supply0 signed abc,ABC;
endmodule
//author : andreib
module input_declaration79( abc,ABC ); input supply0 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration80( abc,ABC ); input supply0 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration81( abc,ABC ); input supply0 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration82( abc,ABC ); input supply0 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration83( abc,ABC ); input supply0 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration84( abc,ABC ); input supply0 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration85( abc,ABC ); input supply0 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration86( abc,ABC ); input supply0 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration87( abc,ABC ); input supply0 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration88( abc,ABC ); input supply0 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration89( abc,ABC ); input supply0 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration90( abc,ABC ); input supply0 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration91( abc,ABC ); input supply0 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration92( abc,ABC ); input supply0 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration93( abc,ABC ); input supply0 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration94( abc,ABC ); input supply0 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration95( abc,ABC ); input supply0 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration96( abc,ABC ); input supply0 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration97( abc,ABC ); input supply0 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration98( abc,ABC ); input supply0 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration99( abc,ABC ); input supply0 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration100( abc,ABC ); input supply0 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration101( abc,ABC ); input supply0 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration102( abc,ABC ); input supply0 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration103( abc,ABC ); input supply0 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration104( abc,ABC ); input supply1 abc,ABC;
endmodule
//author : andreib
module input_declaration105( abc,ABC ); input supply1 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration106( abc,ABC ); input supply1 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration107( abc,ABC ); input supply1 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration108( abc,ABC ); input supply1 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration109( abc,ABC ); input supply1 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration110( abc,ABC ); input supply1 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration111( abc,ABC ); input supply1 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration112( abc,ABC ); input supply1 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration113( abc,ABC ); input supply1 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration114( abc,ABC ); input supply1 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration115( abc,ABC ); input supply1 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration116( abc,ABC ); input supply1 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration117( abc,ABC ); input supply1 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration118( abc,ABC ); input supply1 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration119( abc,ABC ); input supply1 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration120( abc,ABC ); input supply1 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration121( abc,ABC ); input supply1 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration122( abc,ABC ); input supply1 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration123( abc,ABC ); input supply1 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration124( abc,ABC ); input supply1 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration125( abc,ABC ); input supply1 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration126( abc,ABC ); input supply1 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration127( abc,ABC ); input supply1 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration128( abc,ABC ); input supply1 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration129( abc,ABC ); input supply1 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration130( abc,ABC ); input supply1 signed abc,ABC;
endmodule
//author : andreib
module input_declaration131( abc,ABC ); input supply1 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration132( abc,ABC ); input supply1 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration133( abc,ABC ); input supply1 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration134( abc,ABC ); input supply1 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration135( abc,ABC ); input supply1 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration136( abc,ABC ); input supply1 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration137( abc,ABC ); input supply1 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration138( abc,ABC ); input supply1 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration139( abc,ABC ); input supply1 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration140( abc,ABC ); input supply1 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration141( abc,ABC ); input supply1 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration142( abc,ABC ); input supply1 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration143( abc,ABC ); input supply1 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration144( abc,ABC ); input supply1 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration145( abc,ABC ); input supply1 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration146( abc,ABC ); input supply1 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration147( abc,ABC ); input supply1 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration148( abc,ABC ); input supply1 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration149( abc,ABC ); input supply1 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration150( abc,ABC ); input supply1 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration151( abc,ABC ); input supply1 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration152( abc,ABC ); input supply1 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration153( abc,ABC ); input supply1 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration154( abc,ABC ); input supply1 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration155( abc,ABC ); input supply1 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration156( abc,ABC ); input tri abc,ABC;
endmodule
//author : andreib
module input_declaration157( abc,ABC ); input tri [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration158( abc,ABC ); input tri [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration159( abc,ABC ); input tri [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration160( abc,ABC ); input tri [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration161( abc,ABC ); input tri [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration162( abc,ABC ); input tri [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration163( abc,ABC ); input tri [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration164( abc,ABC ); input tri [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration165( abc,ABC ); input tri [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration166( abc,ABC ); input tri [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration167( abc,ABC ); input tri [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration168( abc,ABC ); input tri [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration169( abc,ABC ); input tri [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration170( abc,ABC ); input tri [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration171( abc,ABC ); input tri [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration172( abc,ABC ); input tri [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration173( abc,ABC ); input tri [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration174( abc,ABC ); input tri [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration175( abc,ABC ); input tri [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration176( abc,ABC ); input tri [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration177( abc,ABC ); input tri [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration178( abc,ABC ); input tri [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration179( abc,ABC ); input tri [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration180( abc,ABC ); input tri [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration181( abc,ABC ); input tri [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration182( abc,ABC ); input tri signed abc,ABC;
endmodule
//author : andreib
module input_declaration183( abc,ABC ); input tri signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration184( abc,ABC ); input tri signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration185( abc,ABC ); input tri signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration186( abc,ABC ); input tri signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration187( abc,ABC ); input tri signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration188( abc,ABC ); input tri signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration189( abc,ABC ); input tri signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration190( abc,ABC ); input tri signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration191( abc,ABC ); input tri signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration192( abc,ABC ); input tri signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration193( abc,ABC ); input tri signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration194( abc,ABC ); input tri signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration195( abc,ABC ); input tri signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration196( abc,ABC ); input tri signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration197( abc,ABC ); input tri signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration198( abc,ABC ); input tri signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration199( abc,ABC ); input tri signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration200( abc,ABC ); input tri signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration201( abc,ABC ); input tri signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration202( abc,ABC ); input tri signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration203( abc,ABC ); input tri signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration204( abc,ABC ); input tri signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration205( abc,ABC ); input tri signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration206( abc,ABC ); input tri signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration207( abc,ABC ); input tri signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration208( abc,ABC ); input triand abc,ABC;
endmodule
//author : andreib
module input_declaration209( abc,ABC ); input triand [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration210( abc,ABC ); input triand [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration211( abc,ABC ); input triand [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration212( abc,ABC ); input triand [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration213( abc,ABC ); input triand [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration214( abc,ABC ); input triand [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration215( abc,ABC ); input triand [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration216( abc,ABC ); input triand [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration217( abc,ABC ); input triand [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration218( abc,ABC ); input triand [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration219( abc,ABC ); input triand [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration220( abc,ABC ); input triand [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration221( abc,ABC ); input triand [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration222( abc,ABC ); input triand [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration223( abc,ABC ); input triand [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration224( abc,ABC ); input triand [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration225( abc,ABC ); input triand [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration226( abc,ABC ); input triand [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration227( abc,ABC ); input triand [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration228( abc,ABC ); input triand [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration229( abc,ABC ); input triand [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration230( abc,ABC ); input triand [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration231( abc,ABC ); input triand [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration232( abc,ABC ); input triand [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration233( abc,ABC ); input triand [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration234( abc,ABC ); input triand signed abc,ABC;
endmodule
//author : andreib
module input_declaration235( abc,ABC ); input triand signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration236( abc,ABC ); input triand signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration237( abc,ABC ); input triand signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration238( abc,ABC ); input triand signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration239( abc,ABC ); input triand signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration240( abc,ABC ); input triand signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration241( abc,ABC ); input triand signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration242( abc,ABC ); input triand signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration243( abc,ABC ); input triand signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration244( abc,ABC ); input triand signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration245( abc,ABC ); input triand signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration246( abc,ABC ); input triand signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration247( abc,ABC ); input triand signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration248( abc,ABC ); input triand signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration249( abc,ABC ); input triand signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration250( abc,ABC ); input triand signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration251( abc,ABC ); input triand signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration252( abc,ABC ); input triand signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration253( abc,ABC ); input triand signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration254( abc,ABC ); input triand signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration255( abc,ABC ); input triand signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration256( abc,ABC ); input triand signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration257( abc,ABC ); input triand signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration258( abc,ABC ); input triand signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration259( abc,ABC ); input triand signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration260( abc,ABC ); input trior abc,ABC;
endmodule
//author : andreib
module input_declaration261( abc,ABC ); input trior [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration262( abc,ABC ); input trior [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration263( abc,ABC ); input trior [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration264( abc,ABC ); input trior [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration265( abc,ABC ); input trior [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration266( abc,ABC ); input trior [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration267( abc,ABC ); input trior [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration268( abc,ABC ); input trior [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration269( abc,ABC ); input trior [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration270( abc,ABC ); input trior [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration271( abc,ABC ); input trior [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration272( abc,ABC ); input trior [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration273( abc,ABC ); input trior [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration274( abc,ABC ); input trior [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration275( abc,ABC ); input trior [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration276( abc,ABC ); input trior [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration277( abc,ABC ); input trior [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration278( abc,ABC ); input trior [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration279( abc,ABC ); input trior [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration280( abc,ABC ); input trior [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration281( abc,ABC ); input trior [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration282( abc,ABC ); input trior [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration283( abc,ABC ); input trior [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration284( abc,ABC ); input trior [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration285( abc,ABC ); input trior [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration286( abc,ABC ); input trior signed abc,ABC;
endmodule
//author : andreib
module input_declaration287( abc,ABC ); input trior signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration288( abc,ABC ); input trior signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration289( abc,ABC ); input trior signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration290( abc,ABC ); input trior signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration291( abc,ABC ); input trior signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration292( abc,ABC ); input trior signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration293( abc,ABC ); input trior signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration294( abc,ABC ); input trior signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration295( abc,ABC ); input trior signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration296( abc,ABC ); input trior signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration297( abc,ABC ); input trior signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration298( abc,ABC ); input trior signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration299( abc,ABC ); input trior signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration300( abc,ABC ); input trior signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration301( abc,ABC ); input trior signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration302( abc,ABC ); input trior signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration303( abc,ABC ); input trior signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration304( abc,ABC ); input trior signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration305( abc,ABC ); input trior signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration306( abc,ABC ); input trior signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration307( abc,ABC ); input trior signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration308( abc,ABC ); input trior signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration309( abc,ABC ); input trior signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration310( abc,ABC ); input trior signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration311( abc,ABC ); input trior signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration312( abc,ABC ); input tri0 abc,ABC;
endmodule
//author : andreib
module input_declaration313( abc,ABC ); input tri0 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration314( abc,ABC ); input tri0 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration315( abc,ABC ); input tri0 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration316( abc,ABC ); input tri0 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration317( abc,ABC ); input tri0 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration318( abc,ABC ); input tri0 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration319( abc,ABC ); input tri0 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration320( abc,ABC ); input tri0 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration321( abc,ABC ); input tri0 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration322( abc,ABC ); input tri0 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration323( abc,ABC ); input tri0 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration324( abc,ABC ); input tri0 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration325( abc,ABC ); input tri0 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration326( abc,ABC ); input tri0 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration327( abc,ABC ); input tri0 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration328( abc,ABC ); input tri0 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration329( abc,ABC ); input tri0 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration330( abc,ABC ); input tri0 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration331( abc,ABC ); input tri0 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration332( abc,ABC ); input tri0 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration333( abc,ABC ); input tri0 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration334( abc,ABC ); input tri0 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration335( abc,ABC ); input tri0 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration336( abc,ABC ); input tri0 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration337( abc,ABC ); input tri0 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration338( abc,ABC ); input tri0 signed abc,ABC;
endmodule
//author : andreib
module input_declaration339( abc,ABC ); input tri0 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration340( abc,ABC ); input tri0 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration341( abc,ABC ); input tri0 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration342( abc,ABC ); input tri0 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration343( abc,ABC ); input tri0 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration344( abc,ABC ); input tri0 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration345( abc,ABC ); input tri0 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration346( abc,ABC ); input tri0 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration347( abc,ABC ); input tri0 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration348( abc,ABC ); input tri0 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration349( abc,ABC ); input tri0 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration350( abc,ABC ); input tri0 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration351( abc,ABC ); input tri0 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration352( abc,ABC ); input tri0 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration353( abc,ABC ); input tri0 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration354( abc,ABC ); input tri0 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration355( abc,ABC ); input tri0 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration356( abc,ABC ); input tri0 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration357( abc,ABC ); input tri0 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration358( abc,ABC ); input tri0 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration359( abc,ABC ); input tri0 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration360( abc,ABC ); input tri0 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration361( abc,ABC ); input tri0 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration362( abc,ABC ); input tri0 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration363( abc,ABC ); input tri0 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration364( abc,ABC ); input tri1 abc,ABC;
endmodule
//author : andreib
module input_declaration365( abc,ABC ); input tri1 [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration366( abc,ABC ); input tri1 [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration367( abc,ABC ); input tri1 [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration368( abc,ABC ); input tri1 [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration369( abc,ABC ); input tri1 [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration370( abc,ABC ); input tri1 [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration371( abc,ABC ); input tri1 [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration372( abc,ABC ); input tri1 [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration373( abc,ABC ); input tri1 [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration374( abc,ABC ); input tri1 [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration375( abc,ABC ); input tri1 [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration376( abc,ABC ); input tri1 [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration377( abc,ABC ); input tri1 [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration378( abc,ABC ); input tri1 [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration379( abc,ABC ); input tri1 [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration380( abc,ABC ); input tri1 [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration381( abc,ABC ); input tri1 [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration382( abc,ABC ); input tri1 [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration383( abc,ABC ); input tri1 [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration384( abc,ABC ); input tri1 [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration385( abc,ABC ); input tri1 [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration386( abc,ABC ); input tri1 [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration387( abc,ABC ); input tri1 [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration388( abc,ABC ); input tri1 [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration389( abc,ABC ); input tri1 [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration390( abc,ABC ); input tri1 signed abc,ABC;
endmodule
//author : andreib
module input_declaration391( abc,ABC ); input tri1 signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration392( abc,ABC ); input tri1 signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration393( abc,ABC ); input tri1 signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration394( abc,ABC ); input tri1 signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration395( abc,ABC ); input tri1 signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration396( abc,ABC ); input tri1 signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration397( abc,ABC ); input tri1 signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration398( abc,ABC ); input tri1 signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration399( abc,ABC ); input tri1 signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration400( abc,ABC ); input tri1 signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration401( abc,ABC ); input tri1 signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration402( abc,ABC ); input tri1 signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration403( abc,ABC ); input tri1 signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration404( abc,ABC ); input tri1 signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration405( abc,ABC ); input tri1 signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration406( abc,ABC ); input tri1 signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration407( abc,ABC ); input tri1 signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration408( abc,ABC ); input tri1 signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration409( abc,ABC ); input tri1 signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration410( abc,ABC ); input tri1 signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration411( abc,ABC ); input tri1 signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration412( abc,ABC ); input tri1 signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration413( abc,ABC ); input tri1 signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration414( abc,ABC ); input tri1 signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration415( abc,ABC ); input tri1 signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration416( abc,ABC ); input wire abc,ABC;
endmodule
//author : andreib
module input_declaration417( abc,ABC ); input wire [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration418( abc,ABC ); input wire [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration419( abc,ABC ); input wire [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration420( abc,ABC ); input wire [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration421( abc,ABC ); input wire [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration422( abc,ABC ); input wire [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration423( abc,ABC ); input wire [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration424( abc,ABC ); input wire [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration425( abc,ABC ); input wire [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration426( abc,ABC ); input wire [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration427( abc,ABC ); input wire [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration428( abc,ABC ); input wire [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration429( abc,ABC ); input wire [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration430( abc,ABC ); input wire [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration431( abc,ABC ); input wire [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration432( abc,ABC ); input wire [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration433( abc,ABC ); input wire [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration434( abc,ABC ); input wire [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration435( abc,ABC ); input wire [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration436( abc,ABC ); input wire [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration437( abc,ABC ); input wire [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration438( abc,ABC ); input wire [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration439( abc,ABC ); input wire [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration440( abc,ABC ); input wire [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration441( abc,ABC ); input wire [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration442( abc,ABC ); input wire signed abc,ABC;
endmodule
//author : andreib
module input_declaration443( abc,ABC ); input wire signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration444( abc,ABC ); input wire signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration445( abc,ABC ); input wire signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration446( abc,ABC ); input wire signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration447( abc,ABC ); input wire signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration448( abc,ABC ); input wire signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration449( abc,ABC ); input wire signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration450( abc,ABC ); input wire signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration451( abc,ABC ); input wire signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration452( abc,ABC ); input wire signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration453( abc,ABC ); input wire signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration454( abc,ABC ); input wire signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration455( abc,ABC ); input wire signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration456( abc,ABC ); input wire signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration457( abc,ABC ); input wire signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration458( abc,ABC ); input wire signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration459( abc,ABC ); input wire signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration460( abc,ABC ); input wire signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration461( abc,ABC ); input wire signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration462( abc,ABC ); input wire signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration463( abc,ABC ); input wire signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration464( abc,ABC ); input wire signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration465( abc,ABC ); input wire signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration466( abc,ABC ); input wire signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration467( abc,ABC ); input wire signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration468( abc,ABC ); input wand abc,ABC;
endmodule
//author : andreib
module input_declaration469( abc,ABC ); input wand [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration470( abc,ABC ); input wand [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration471( abc,ABC ); input wand [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration472( abc,ABC ); input wand [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration473( abc,ABC ); input wand [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration474( abc,ABC ); input wand [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration475( abc,ABC ); input wand [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration476( abc,ABC ); input wand [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration477( abc,ABC ); input wand [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration478( abc,ABC ); input wand [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration479( abc,ABC ); input wand [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration480( abc,ABC ); input wand [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration481( abc,ABC ); input wand [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration482( abc,ABC ); input wand [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration483( abc,ABC ); input wand [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration484( abc,ABC ); input wand [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration485( abc,ABC ); input wand [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration486( abc,ABC ); input wand [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration487( abc,ABC ); input wand [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration488( abc,ABC ); input wand [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration489( abc,ABC ); input wand [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration490( abc,ABC ); input wand [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration491( abc,ABC ); input wand [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration492( abc,ABC ); input wand [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration493( abc,ABC ); input wand [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration494( abc,ABC ); input wand signed abc,ABC;
endmodule
//author : andreib
module input_declaration495( abc,ABC ); input wand signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration496( abc,ABC ); input wand signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration497( abc,ABC ); input wand signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration498( abc,ABC ); input wand signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration499( abc,ABC ); input wand signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration500( abc,ABC ); input wand signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration501( abc,ABC ); input wand signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration502( abc,ABC ); input wand signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration503( abc,ABC ); input wand signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration504( abc,ABC ); input wand signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration505( abc,ABC ); input wand signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration506( abc,ABC ); input wand signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration507( abc,ABC ); input wand signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration508( abc,ABC ); input wand signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration509( abc,ABC ); input wand signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration510( abc,ABC ); input wand signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration511( abc,ABC ); input wand signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration512( abc,ABC ); input wand signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration513( abc,ABC ); input wand signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration514( abc,ABC ); input wand signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration515( abc,ABC ); input wand signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration516( abc,ABC ); input wand signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration517( abc,ABC ); input wand signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration518( abc,ABC ); input wand signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration519( abc,ABC ); input wand signed [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration520( abc,ABC ); input wor abc,ABC;
endmodule
//author : andreib
module input_declaration521( abc,ABC ); input wor [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration522( abc,ABC ); input wor [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration523( abc,ABC ); input wor [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration524( abc,ABC ); input wor [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration525( abc,ABC ); input wor [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration526( abc,ABC ); input wor [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration527( abc,ABC ); input wor [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration528( abc,ABC ); input wor [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration529( abc,ABC ); input wor [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration530( abc,ABC ); input wor [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration531( abc,ABC ); input wor [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration532( abc,ABC ); input wor [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration533( abc,ABC ); input wor [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration534( abc,ABC ); input wor [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration535( abc,ABC ); input wor [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration536( abc,ABC ); input wor [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration537( abc,ABC ); input wor [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration538( abc,ABC ); input wor [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration539( abc,ABC ); input wor [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration540( abc,ABC ); input wor [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration541( abc,ABC ); input wor [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration542( abc,ABC ); input wor [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration543( abc,ABC ); input wor [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration544( abc,ABC ); input wor [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration545( abc,ABC ); input wor [ "str" : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration546( abc,ABC ); input wor signed abc,ABC;
endmodule
//author : andreib
module input_declaration547( abc,ABC ); input wor signed [ 2 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration548( abc,ABC ); input wor signed [ 2 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration549( abc,ABC ); input wor signed [ 2 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration550( abc,ABC ); input wor signed [ 2 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration551( abc,ABC ); input wor signed [ 2 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration552( abc,ABC ); input wor signed [ +3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration553( abc,ABC ); input wor signed [ +3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration554( abc,ABC ); input wor signed [ +3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration555( abc,ABC ); input wor signed [ +3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration556( abc,ABC ); input wor signed [ +3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration557( abc,ABC ); input wor signed [ 2-1 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration558( abc,ABC ); input wor signed [ 2-1 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration559( abc,ABC ); input wor signed [ 2-1 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration560( abc,ABC ); input wor signed [ 2-1 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration561( abc,ABC ); input wor signed [ 2-1 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration562( abc,ABC ); input wor signed [ 1?2:3 : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration563( abc,ABC ); input wor signed [ 1?2:3 : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration564( abc,ABC ); input wor signed [ 1?2:3 : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration565( abc,ABC ); input wor signed [ 1?2:3 : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration566( abc,ABC ); input wor signed [ 1?2:3 : "str" ] abc,ABC;
endmodule
//author : andreib
module input_declaration567( abc,ABC ); input wor signed [ "str" : 1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration568( abc,ABC ); input wor signed [ "str" : +1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration569( abc,ABC ); input wor signed [ "str" : 2-1 ] abc,ABC;
endmodule
//author : andreib
module input_declaration570( abc,ABC ); input wor signed [ "str" : 1?2:3 ] abc,ABC;
endmodule
//author : andreib
module input_declaration571( abc,ABC ); input wor signed [ "str" : "str" ] abc,ABC;
endmodule
