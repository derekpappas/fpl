`include "a.vh"

module a ();
wire a = `A;
endmodule