// Test type: case_statement - casez - expression:null
// Vparser rule name:
// Author: andreib
module case_statement41;
reg a;
initial casez(a)
	4'bzZ?0:;
	endcase
endmodule
