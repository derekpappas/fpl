`include "defines.v"

module n1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 262
  output [1 - 1:0] ar_sa0_s10;
  m1 m10(.ar_sa0_s10(ar_sa0_s10));
  `include "n1.logic.vh"
endmodule

