`define A 1'b1