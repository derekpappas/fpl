//test type : number binary_operator_** number
//vparser rule name : 
//author : Bogdan Mereghea
module binary_operator37;
    reg a;
    initial begin 
        a = 1'b1 ** 1'd2; 
    end
endmodule
