//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : ddr_ctrl.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module ddr_ctrl(dc_dbcdummy5,
                dc_dbdummy5);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 31
  output dc_dbcdummy5;
  output dc_dbdummy5;
  `include "ddr_ctrl.logic.v"
endmodule

