// Test type: Continuous assignment - pl1, wk0 - list_of_net_assignments - 2 elements
// Vparser rule name:
// Author: andreib
module continuous422;
wire a,b;
assign (pull1, weak0) a=1'b1, b=1'b0;
endmodule
