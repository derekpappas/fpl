a.vhd
b.vhd
c.vhd
top.vhd
