`define outside
module
if( 
`define inside 24
`inside > 10);
endmodule
`undef outside
`undef inside
