// Test type: Strings - 2 chars String
// Vparser rule name:
// Author: andreib
module stringtest;
reg [8*32:1] stringvar;
initial begin
stringvar = "az";
end
endmodule
