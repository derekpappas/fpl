// Test type: Binary Numbers - signed number base lower case
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=3'sb101;
endmodule
