module x;
`default_nettype
endmodule
