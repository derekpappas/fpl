// Test type: Decimal Numbers - Decimal number with underscores
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=48_3_;
endmodule
