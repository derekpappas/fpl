`include "defines.v"

module m_im();
// Location of source csl unit: file name = mbist_datapath.csl line number = 76
// The depth of memory module m_im is of illegal type. Depth set to 1.
// The width of memory module m_im is of illegal type. Width set to 1.
  endmodule

