// Test type: blocking_assignment - delay control - expression
// Vparser rule name:
// Author: andreib
module blocking_assignment2;
reg a;
initial a=#10 2;
endmodule
