module testbench_gate_instantiation;
    gate_instantiation0 gate_instantiation_instance0();
    gate_instantiation1 gate_instantiation_instance1();
    gate_instantiation2 gate_instantiation_instance2();
    gate_instantiation3 gate_instantiation_instance3();
    gate_instantiation4 gate_instantiation_instance4();
    gate_instantiation5 gate_instantiation_instance5();
    gate_instantiation6 gate_instantiation_instance6();
    gate_instantiation7 gate_instantiation_instance7();
    gate_instantiation8 gate_instantiation_instance8();
    gate_instantiation9 gate_instantiation_instance9();
    gate_instantiation10 gate_instantiation_instance10();
    gate_instantiation11 gate_instantiation_instance11();
    gate_instantiation12 gate_instantiation_instance12();
    gate_instantiation13 gate_instantiation_instance13();
    gate_instantiation14 gate_instantiation_instance14();
    gate_instantiation15 gate_instantiation_instance15();
    gate_instantiation16 gate_instantiation_instance16();
    gate_instantiation17 gate_instantiation_instance17();
    gate_instantiation18 gate_instantiation_instance18();
    gate_instantiation19 gate_instantiation_instance19();
    gate_instantiation20 gate_instantiation_instance20();
    gate_instantiation21 gate_instantiation_instance21();
    gate_instantiation22 gate_instantiation_instance22();
    gate_instantiation23 gate_instantiation_instance23();
    gate_instantiation24 gate_instantiation_instance24();
    gate_instantiation25 gate_instantiation_instance25();
    gate_instantiation26 gate_instantiation_instance26();
    gate_instantiation27 gate_instantiation_instance27();
    gate_instantiation28 gate_instantiation_instance28();
    gate_instantiation29 gate_instantiation_instance29();
    gate_instantiation30 gate_instantiation_instance30();
    gate_instantiation31 gate_instantiation_instance31();
    gate_instantiation32 gate_instantiation_instance32();
    gate_instantiation33 gate_instantiation_instance33();
    gate_instantiation34 gate_instantiation_instance34();
    gate_instantiation35 gate_instantiation_instance35();
    gate_instantiation36 gate_instantiation_instance36();
    gate_instantiation37 gate_instantiation_instance37();
    gate_instantiation38 gate_instantiation_instance38();
    gate_instantiation39 gate_instantiation_instance39();
endmodule
//@
//author : andreib
module gate_instantiation0(a,b);
parameter id_a=1;
inout a,b;
tranif0 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation1(a,b);
parameter id_a=1;
inout a,b;
tranif0 # 2 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation2(a,b);
parameter id_a=1;
inout a,b;
tranif0 # 1.2e1 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation3(a,b);
parameter id_a=1;
inout a,b;
tranif0 # id_a ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation4(a,b);
parameter id_a=1;
inout a,b;
tranif0 #( 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation5(a,b);
parameter id_a=1;
inout a,b;
tranif0 #( 1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation6(a,b);
parameter id_a=1;
inout a,b;
tranif0 #( 1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation7(a,b);
parameter id_a=1;
inout a,b;
tranif0 #( 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation8(a,b);
parameter id_a=1;
inout a,b;
tranif0 #( 1 : +1 : 2+1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation9(a,b);
parameter id_a=1;
inout a,b;
tranif0 #( 1 : +1 : 2+1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation10(a,b);
parameter id_a=1;
inout a,b;
tranif1 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation11(a,b);
parameter id_a=1;
inout a,b;
tranif1 # 2 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation12(a,b);
parameter id_a=1;
inout a,b;
tranif1 # 1.2e1 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation13(a,b);
parameter id_a=1;
inout a,b;
tranif1 # id_a ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation14(a,b);
parameter id_a=1;
inout a,b;
tranif1 #( 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation15(a,b);
parameter id_a=1;
inout a,b;
tranif1 #( 1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation16(a,b);
parameter id_a=1;
inout a,b;
tranif1 #( 1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation17(a,b);
parameter id_a=1;
inout a,b;
tranif1 #( 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation18(a,b);
parameter id_a=1;
inout a,b;
tranif1 #( 1 : +1 : 2+1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation19(a,b);
parameter id_a=1;
inout a,b;
tranif1 #( 1 : +1 : 2+1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation20(a,b);
parameter id_a=1;
inout a,b;
rtranif1 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation21(a,b);
parameter id_a=1;
inout a,b;
rtranif1 # 2 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation22(a,b);
parameter id_a=1;
inout a,b;
rtranif1 # 1.2e1 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation23(a,b);
parameter id_a=1;
inout a,b;
rtranif1 # id_a ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation24(a,b);
parameter id_a=1;
inout a,b;
rtranif1 #( 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation25(a,b);
parameter id_a=1;
inout a,b;
rtranif1 #( 1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation26(a,b);
parameter id_a=1;
inout a,b;
rtranif1 #( 1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation27(a,b);
parameter id_a=1;
inout a,b;
rtranif1 #( 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation28(a,b);
parameter id_a=1;
inout a,b;
rtranif1 #( 1 : +1 : 2+1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation29(a,b);
parameter id_a=1;
inout a,b;
rtranif1 #( 1 : +1 : 2+1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation30(a,b);
parameter id_a=1;
inout a,b;
rtranif0 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation31(a,b);
parameter id_a=1;
inout a,b;
rtranif0 # 2 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation32(a,b);
parameter id_a=1;
inout a,b;
rtranif0 # 1.2e1 ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation33(a,b);
parameter id_a=1;
inout a,b;
rtranif0 # id_a ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation34(a,b);
parameter id_a=1;
inout a,b;
rtranif0 #( 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation35(a,b);
parameter id_a=1;
inout a,b;
rtranif0 #( 1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation36(a,b);
parameter id_a=1;
inout a,b;
rtranif0 #( 1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation37(a,b);
parameter id_a=1;
inout a,b;
rtranif0 #( 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation38(a,b);
parameter id_a=1;
inout a,b;
rtranif0 #( 1 : +1 : 2+1 , 1 ) ( a , b , 1'b1 );
endmodule
//author : andreib
module gate_instantiation39(a,b);
parameter id_a=1;
inout a,b;
rtranif0 #( 1 : +1 : 2+1 , 1 : +1 : 2+1 ) ( a , b , 1'b1 );
endmodule
