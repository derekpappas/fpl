// Test type: Decimal Numbers - signed decimal number  
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'sd16;
endmodule
