`define a \`include
module `a;
//reg x;
endmodule

