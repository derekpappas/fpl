// Test type: case_statement - casez - 2 x expression:null
// Vparser rule name:
// Author: andreib
module case_statement51;
reg a;
initial casez(a)
	4'bzZ?0:;
	4'b0001:;
	endcase
endmodule
