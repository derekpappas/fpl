// Test type: Expression - string
// Vparser rule name:
// Author: andreib
module expressiontest;
reg [8*31:0] string;
initial begin
string = "This is a string";
end
endmodule
