`define x mememumu
module \A ;
`x
endmodule
