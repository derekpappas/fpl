// Test type: Binary Numbers - Size specified
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=8'b10110110;
endmodule
