//test type : module_declaration
//vparser rule name : 
//author : Codrin
(* a *)
(* a = 1 *)
(* a, b *)
module declaration_020;
endmodule
