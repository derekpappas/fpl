// Test type: Continuous assignment - 1 mintypmax - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous7;
wire a;
assign #(1) a=1'b1;
endmodule
