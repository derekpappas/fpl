// Test type: delay_control - (mintypmax) - expression
// Vparser rule name:
// Author: andreib
module delay_control4;
reg a;
initial #(1) a=1'b1;
endmodule
