`define identifier xx
module x`identifier;
reg a,b;
wire c;
and #1 (a,b,c);
endmodule
