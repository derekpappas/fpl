`include "defines.v"

module p1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 274
  output [1 - 1:0] ar_sa0_s10;
  o1 o10(.ar_sa0_s10(ar_sa0_s10));
  `include "p1.logic.vh"
endmodule

