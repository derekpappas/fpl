//test type : {constant_expression}
//vparser rule name : 
//author : Bogdan Mereghea
module constant_concatenation1;
    wire a;
    assign a = {1'b1};
endmodule
