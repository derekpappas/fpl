-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./msi_rx_cslc_generated/code/vhdl/sfd_trans.vhd
-- FILE GENERATED ON : Thu Jun 19 15:32:42 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \sfd_trans\ is
  port(\lbdummy3\ : in csl_bit);
begin
end entity;

architecture \sfd_trans_logic\ of \sfd_trans\ is
begin
end architecture;

