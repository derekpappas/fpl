`default_nettype tri
`celldefine
module yyy;
`include "../legal/default_nettype06.v"
wire x;
`celldefine
wire t;
`default_nettype none
endmodule
