//au.vh