// Test type: conditional_statement - if(expr) statement else statement
// Vparser rule name:
// Author: andreib
module conditional_statement6;
reg a,b,c;
initial if(a==b) c=1;
else c=0;
endmodule
