`define number 1
module x;
reg a,b;
wire c;
and #1`number (a,b,c);
endmodule
