// Test type: delay_or_event_control - event_control
// Vparser rule name:
// Author: andreib
module delay_or_event_control3;
reg a,clk;
initial @clk a=1'b1;
endmodule
