`include "defines.v"

module u_b(p_b_in);
// Location of source csl unit: file name = ar3b.csl line number = 34
  input [2 - 1:0] p_b_in;
  `include "u_b.logic.v"
endmodule

