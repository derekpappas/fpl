// Test type: Continuous assignment - list_of_net_assignments - 2 elements
// Vparser rule name:
// Author: andreib
module continuous2;
wire a,b;
assign a=1'b1, b=1'b0;
endmodule
