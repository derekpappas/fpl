//test type : module_or_generate_item ::= module_or_generate_item_declaration (genvar_declaration)
//vparser rule name : 
//author : Codrin
module test_0230;
 (* generated = 1 *)
 genvar i;
endmodule
