// Test type: Octal Numbers - 1 number
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=3'o5;
endmodule
