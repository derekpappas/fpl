-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top_cslc_generated/code/vhdl/uu.vhd
-- FILE GENERATED ON : Sat Mar 14 18:10:30 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \uu\ is
  port(\sel\ : in csl_bit_vector(10#2# - 10#1# downto 10#0#);
       \irc_reset\ : in csl_bit;
       \irc_clock\ : in csl_bit;
       \iin_pinx\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \iin_piny\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \iout_pinx\ : out csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \iout_piny\ : out csl_bit_vector(10#8# - 10#1# downto 10#0#));
begin
end entity;

architecture \uu_logic\ of \uu\ is
begin
end architecture;

