module x;
`line 1 "" 1
endmodule
