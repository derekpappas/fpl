`include "defines.v"

module a0(sa0);
// Location of source csl unit: file name = temp.csl line number = 1
  input sa0;
  `include "a0.logic.vh"
endmodule

