`define x 
`define y \��
module modul;
//reg `x = 1;
reg `y;
endmodule
