//test type : port_declaration
//vparser rule name : 
//author : Codrin
module declaration_0100(x);
 (* a , b, c = 1 *) input x;
endmodule
