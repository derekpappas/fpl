// Test type: Hex Numbers - underscore within value
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8'h1___9;
endmodule
