`include "defines.v"

module w1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 318
  output [1 - 1:0] ar_sa0_s10;
  v1 v10(.ar_sa0_s10(ar_sa0_s10));
  `include "w1.logic.vh"
endmodule

