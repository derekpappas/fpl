//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : spi_cntl_cluster.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module spi_cntl_cluster();
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 16
  spi_cntl spi_cntl();
  spi_cntl_lba spi_cntl_lba();
  msi_fabric_if spi_cntl_fab();
  `include "spi_cntl_cluster.logic.v"
endmodule

