// Test type: Hex Numbers - 2 numbers upper case base
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8'HA3;
endmodule
