//test type : hierarchical_identifier binary_operator_** hierarchical_identifier
//vparser rule name : 
//author : Bogdan Mereghea
module binary_operator12;
    reg a, b, c;
    initial begin 
    a = b ** 1'd2; 
    end
endmodule
