module b(y);
input y;
endmodule
