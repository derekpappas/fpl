module x;
endmodule
`nounconnected_drive
module t;
endmodule
