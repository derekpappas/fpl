`include "defines.v"

module eu();
// Location of source csl unit: file name = /Volumes/s2/unfuddle_ssm_repo/ssm_ssmrepo/ssm/hw/ssm/ssm_demo.csl line number = 91
  `include "eu.logic.vh"
endmodule

