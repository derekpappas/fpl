`define comment /
module x;
reg a,b;
wire c;
/`comment (a,b,c);
endmodule
