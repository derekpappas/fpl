// Test type: Binary Numbers - No size specified upper case base
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a='B1011;
endmodule
