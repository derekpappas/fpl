//test type : module_or_generate_item ::= continuous_assign
//vparser rule name : 
//author : Codrin
module test_0270;
 (* integers = 1 *) wire a;
 assign a = 5'd18;
endmodule
