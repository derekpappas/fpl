`include "b.vh"

module b ();
wire b = `B;
endmodule