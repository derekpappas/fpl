//qm.vh