`include "defines.v"

module k1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 244
  output [1 - 1:0] ar_sa0_s10;
  j1 j10(.ar_sa0_s10(ar_sa0_s10));
  `include "k1.logic.vh"
endmodule

