// Test type: Continuous assignment - st0, sup1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous76;
wire a;
assign (strong0, supply1) a=1'b1;
endmodule
