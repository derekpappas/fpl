//test type : module_or_generate_item ::= module_or_generate_item_declaration (reg_declaration)
//vparser rule name : 
//author : Codrin
module test_0160;
 (* fsm_state=1 *) reg [3:0] state2, state3;
endmodule
