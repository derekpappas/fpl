// Test type: procedural continuous assignment - assign variable assignment
// Vparser rule name:
// Author: andreib
module procedural_continuous_assignment1;
reg a;
initial assign a=1'b1;
endmodule
