`celldefine
module xxx;
endmodule
`include "../legal/celldef19.v"
`celldefine
`include "../legal/celldef19.v"
`celldefine
`include "../legal/celldef19.v"
`celldefine
`include "../legal/celldef19.v"
`celldefine
`include "../legal/celldef19.v"
module yyy;
endmodule
`resetall
