// Test type: Continuous assignment - sup0, pl1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous46;
wire a;
assign (supply0, pull1) a=1'b1;
endmodule
