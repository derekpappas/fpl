r_pc.vhd
m_im.vhd
rf.vhd
rf_register_file_memory.vhd
u_arith.vhd
u_logic.vhd
u_mux41.vhd
u_cmp.vhd
u_sh.vhd
u_alu_sh_cmp.vhd
u_control.vhd
u_mbist.vhd
