// Test type: Decimal Numbers - space between size and base
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=32 'd16;
endmodule
