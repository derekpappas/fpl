// Test type: Hex Numbers - ? and z digit
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=16'h9z?Z;
endmodule
