`include "defines.v"

module q0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 113
  input [1 - 1:0] ar_sa0_s10;
  p0 p0(.ar_sa0_s10(ar_sa0_s10));
  `include "q0.logic.vh"
endmodule

