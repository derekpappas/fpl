`include "defines.v"

module u3();
// Location of source csl unit: file name = ar16.csl line number = 43
  `include "u3.logic.v"
endmodule

