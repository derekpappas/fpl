// Test type: Decimal Numbers - Large decimal number
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=1234567890;
endmodule
