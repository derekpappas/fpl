// Test type: net_assignment - primary
// Vparser rule name:
// Author: andreib
module netasign1;
wire a;
assign a=2;
endmodule
