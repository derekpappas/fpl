//test type : specify_block_declaration
//author : Dramba Doru-Gabriel
module setuphold_timing_check0(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" );endspecify
endmodule
module setuphold_timing_check1(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , );endspecify
endmodule
module setuphold_timing_check2(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , );endspecify
endmodule
module setuphold_timing_check3(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , );endspecify
endmodule
module setuphold_timing_check4(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , );endspecify
endmodule
module setuphold_timing_check5(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , , );endspecify
endmodule
module setuphold_timing_check6(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check7(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check8(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check9(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check10(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check11(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check12(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check13(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check14(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check15(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check16(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 );endspecify
endmodule
module setuphold_timing_check17(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , );endspecify
endmodule
module setuphold_timing_check18(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , , );endspecify
endmodule
module setuphold_timing_check19(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check20(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check21(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check22(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check23(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check24(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check25(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check26(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check27(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check28(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check29(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 );endspecify
endmodule
module setuphold_timing_check30(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , );endspecify
endmodule
module setuphold_timing_check31(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , );endspecify
endmodule
module setuphold_timing_check32(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , , );endspecify
endmodule
module setuphold_timing_check33(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check34(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check35(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check36(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check37(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check38(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check39(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check40(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check41(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check42(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check43(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 );endspecify
endmodule
module setuphold_timing_check44(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , );endspecify
endmodule
module setuphold_timing_check45(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , , );endspecify
endmodule
module setuphold_timing_check46(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check47(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check48(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check49(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check50(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check51(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check52(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check53(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check54(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check55(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check56(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check57(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check58(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , );endspecify
endmodule
module setuphold_timing_check59(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , );endspecify
endmodule
module setuphold_timing_check60(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , , );endspecify
endmodule
module setuphold_timing_check61(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check62(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check63(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check64(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check65(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check66(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check67(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check68(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check69(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check70(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check71(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 );endspecify
endmodule
module setuphold_timing_check72(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , );endspecify
endmodule
module setuphold_timing_check73(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , , );endspecify
endmodule
module setuphold_timing_check74(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check75(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check76(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check77(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check78(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check79(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check80(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check81(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check82(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check83(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check84(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 );endspecify
endmodule
module setuphold_timing_check85(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , );endspecify
endmodule
module setuphold_timing_check86(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , );endspecify
endmodule
module setuphold_timing_check87(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , , );endspecify
endmodule
module setuphold_timing_check88(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check89(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check90(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check91(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check92(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check93(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check94(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check95(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check96(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check97(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check98(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 );endspecify
endmodule
module setuphold_timing_check99(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , );endspecify
endmodule
module setuphold_timing_check100(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , , );endspecify
endmodule
module setuphold_timing_check101(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check102(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check103(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check104(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier , );endspecify
endmodule
module setuphold_timing_check105(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check106(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier , inoutPortIdentifier[2:2:2] );endspecify
endmodule
module setuphold_timing_check107(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] );endspecify
endmodule
module setuphold_timing_check108(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , );endspecify
endmodule
module setuphold_timing_check109(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier );endspecify
endmodule
module setuphold_timing_check110(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  reg ter;
  specify $setuphold( inoutPortIdentifier , inoutPortIdentifier , "timing=expression" , "timing=expression" , inoutPortIdentifier , 3:3:3 , 2:2:2 , inoutPortIdentifier[3:3:3] , inoutPortIdentifier[2:2:2] );endspecify
endmodule
