// Test type: Binary Numbers - Underscore within size and value
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=1_2'b011_010_000_111;
endmodule
