u_ff.vhd
u_dep.vhd
