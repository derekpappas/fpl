// Test type: Decimal Numbers - size with underscore
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=3__2'd16;
endmodule
