`include "defines.v"

module a(p);
// Location of source csl unit: file name = br_invalid.csl line number = 6
  input [4 - 1:0] p;
  `include "a.logic.v"
endmodule

