`include "defines.v"

module z0();
// Location of source csl unit: file name = temp.csl line number = 341
  wire [1 - 1:0] ar_sa0_s10;
  y0 y0(.ar_sa0_s10(ar_sa0_s10));
  y1 y10(.ar_sa0_s10(ar_sa0_s10));
  `include "z0.logic.vh"
endmodule

