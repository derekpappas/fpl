//test type : task_item_declaration ::= output_declaration
//vparser rule name : 
//author : Codrin
//fixed by: Gabrield
module test_0430;
 task add;
  (* cout, cin *) output sum;
  ;
 endtask
endmodule
