-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./d_cslc_generated/code/vhdl/a.vhd
-- FILE GENERATED ON : Tue Apr 14 20:40:05 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \a\ is
  port(\ck\ : in csl_bit;
       \reset\ : in csl_bit);
begin
end entity;

architecture \a_logic\ of \a\ is
begin
end architecture;

