//test type : module_or_generate_item ::= module_or_generate_item_declaration (time_declaration)
//vparser rule name : 
//author : Codrin
module test_0200;
 (* rtime = 1, treal =0, rinteger = 0 *) time hist[1:100];
endmodule
