`default_nettype tri
module x;
`default_nettype tri0
wire q;
`default_nettype tri1
wire w;
`default_nettype wand
wire e;
`default_nettype triand
wire r;
`default_nettype wor
wire t;
`default_nettype trior
wire y;
`default_nettype trireg
endmodule
