//test type : {expression}
//vparser rule name : 
//author : Bogdan Mereghea
module concatenation1;
    wire a;
    assign a = {1'b1};
endmodule
