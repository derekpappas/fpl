// Test type: Hex Numbers - all numbers
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=4096'h01234567890aAbBcCdDeEfF;
endmodule
