// Test type: Continuous assignment - sup0, st1 - list_of_net_assignments - 3 elements
// Vparser rule name:
// Author: andreib
module continuous33;
wire a,b,c;
assign (supply0, strong1) a=1'b1, b=1'b0, c=1'd2;
endmodule
