`include "defines.v"

module output_cell();
// Location of source csl unit: file name = generated/vizzini_core.csl line number = 162
  `include "output_cell.logic.v"
endmodule

