// Test type: Real numbers - exponent case
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=12.3E12;
endmodule
