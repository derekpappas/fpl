// Test type: always statement - blocking_assignment - no attribute instance
// Vparser rule name:
// Author: andreib
module alwcon1;
reg [7:0]a;
always a=2;
endmodule
