// Test type: Hex Numbers - variations of letter case in signed and base
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8'Sh3F;
endmodule
