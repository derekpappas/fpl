`include "defines.v"

module rfmux();
// Location of source csl unit: file name = IPX2400.csl line number = 66
  `include "rfmux.logic.v"
endmodule

