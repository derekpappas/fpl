// Test type: Decimal Numbers - no size decimal base upper case
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a='D79;
endmodule
