// Test type: Decimal Numbers - upper case signed and decimal base
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'SD2___9;
endmodule
