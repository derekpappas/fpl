//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : spi_cntl.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module spi_cntl(lbadummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 28
  input lbadummy3;
  `include "spi_cntl.logic.v"
endmodule

