//32-bit shifter 
module shifter(sh_out, op, pos, sh_in, clk);
    input [31:0] sh_in;
    input [2:0] op;
    input [4:0] pos;
    input clk;
    output [31:0] sh_out;
    
    always@(clk) begin
            
    end
endmodule