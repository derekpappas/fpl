//test type : non_port_module_item ::= specparam_declaration
//vparser rule name : 
//author : Codrin
//modified by: Gabriel
module test_0390;
// specify
 (* param *)
   specparam min_time = 3;
// endspecify
endmodule
