-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top_cslc_generated/code/vhdl/u23.vhd
-- FILE GENERATED ON : Tue Mar 10 20:48:07 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u23\ is
  port(\ifc_in3_pi1\ : in csl_bit_vector(10#2# - 10#1# downto 10#0#);
       \ifc_in3_pi2\ : in csl_bit_vector(10#4# - 10#1# downto 10#0#);
       \ifc_in3_pi3\ : in csl_bit;
       \ifc_out3_po1\ : out csl_bit_vector(10#2# - 10#1# downto 10#0#);
       \ifc_out3_po2\ : out csl_bit_vector(10#4# - 10#1# downto 10#0#);
       \ifc_out3_po3\ : out csl_bit;
       \ifc_in1_ar_pi1_s1\ : in csl_bit_vector(10#2# - 10#1# downto 10#0#);
       \ifc_in1_ar_pi2_s2\ : in csl_bit_vector(10#4# - 10#1# downto 10#0#);
       \ifc_in1_ar_pi3_s3\ : in csl_bit_vector(10#1# - 10#1# downto 10#0#));
begin
end entity;

architecture \u23_logic\ of \u23\ is

  component \u22\ is
    port(\ifc_in1_ar_pi1_s1\ : in csl_bit_vector(10#2# - 10#1# downto 10#0#);
         \ifc_in1_ar_pi2_s2\ : in csl_bit_vector(10#4# - 10#1# downto 10#0#);
         \ifc_in1_ar_pi3_s3\ : in csl_bit_vector(10#1# - 10#1# downto 10#0#));
  end component;
begin
  -- In file 'TO BE IMPLEMENTED':48 instance name must difer from the instantiated obejct name.
end architecture;

