module a(o);
    wire x;
    output o;
    assign o = b.y;
endmodule
