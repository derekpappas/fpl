`include "defines.v"

module y0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 173
  input [1 - 1:0] ar_sa0_s10;
  x0 x0(.ar_sa0_s10(ar_sa0_s10));
  `include "y0.logic.vh"
endmodule

