// Test type: Octal Numbers - z and ? digit in octal value
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=12'o7z?Z;
endmodule
