//test type : function_port_list ::= input_declaration
//vparser rule name : 
//author : Codrin
module test_0400;
 function [7:0] pow(
  (* width = 8, size *)
  input nr);
  pow = 8'b0;
 endfunction
endmodule
