//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : sd_flash.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module sd_flash(lbdummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 20
  input lbdummy3;
  `include "sd_flash.logic.v"
endmodule

