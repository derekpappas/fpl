`include "defines.v"

module execu();
// Location of source csl unit: file name = IPX2400.csl line number = 34
  `include "execu.logic.v"
endmodule

