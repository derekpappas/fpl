// Test type: Expression - primary - number
// Vparser rule name:
// Author: andreib
module expressiontest;
wire a;
assign a=6'd32;
endmodule
