`unconnected_drive pull1
module x;
endmodule
`nounconnected_drive
module xx;
endmodule
`nounconnected_drive
