// Test type: Hex Numbers - space between base and value
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8'h 3E;
endmodule
