a.vhd
b.vhd
c.vhd
d.vhd
