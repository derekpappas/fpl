`include "defines.v"

module r0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 119
  input [1 - 1:0] ar_sa0_s10;
  q0 q0(.ar_sa0_s10(ar_sa0_s10));
  `include "r0.logic.vh"
endmodule

