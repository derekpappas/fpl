//cl.vh