//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : nios.v
//FILE GENERATED ON : Wed Jul  9 20:26:20 2008

`include "defines.v"

module nios();
// Location of source csl unit: file name = generated/mitch.csl line number = 26
  `include "nios.logic.v"
endmodule

