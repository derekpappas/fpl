//test type : module_or_generate_item ::= module_or_generate_item_declaration (integer_declaration)
//vparser rule name : 
//author : Codrin
module test_0180;
 (* nets = 1 *) wire out;
 assign out = 4'sd21;
endmodule
