// Test type: Continuous assignment - sup0, wk1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous61;
wire a;
assign (supply0, weak1) a=1'b1;
endmodule
