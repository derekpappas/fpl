`include "defines.v"

module u0();
// Location of source csl unit: file name = ar16.csl line number = 31
  `include "u0.logic.v"
endmodule

