--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : a.vh
--FILE GENERATED ON : Wed Jan 20 06:20:06 2010

a.vhd
