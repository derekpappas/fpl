//test type : operator_~^ number
//vparser rule name : 
//author : Bogdan Mereghea
module unary_operator21;
    wire a;
    assign a = ~^1'b1;
endmodule
