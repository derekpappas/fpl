// Test type: Real numbers - simple exponential number
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1e9;
endmodule
