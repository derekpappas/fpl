-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_top_cslc_generated/code/vhdl/u_d.vhd
-- FILE GENERATED ON : Wed Mar 11 20:42:30 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_d\ is
  port(\p_d_in1\ : in csl_bit_vector(10#2# - 10#1# downto 10#0#);
       \p_d_out\ : out csl_bit);
begin
end entity;

architecture \u_d_logic\ of \u_d\ is
begin
end architecture;

