// Test type: Decimal Numbers - x-digit with underscore
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'dx__;
endmodule
