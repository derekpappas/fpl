//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : mfd_sec.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module mfd_sec(lbdummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 10
  input lbdummy3;
  `include "mfd_sec.logic.v"
endmodule

