`include "defines.v"

module input_cell();
// Location of source csl unit: file name = generated/vizzini_core.csl line number = 150
  `include "input_cell.logic.v"
endmodule

