//test type : module_or_generate_item ::= function_call
//vparser rule name : 
//author : Codrin
module test_0320;
 wire a, b, c;
 assign a = add (* mode = "cla" *) (b, c);
endmodule
