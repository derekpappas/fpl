-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_mbist_cslc_generated/code/vhdl/u_es.vhd
-- FILE GENERATED ON : Tue Feb 17 20:24:21 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_es\ is
  port(\p_c\ : in csl_bit_vector(10#7# downto 10#0#);
       \p_ec\ : out csl_bit_vector(10#15# downto 10#0#));
begin
end entity;

architecture \u_es_logic\ of \u_es\ is
begin
end architecture;

