`include "defines.v"

module b1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 189
  output [1 - 1:0] ar_sa0_s10;
  a1 a10(.s10(ar_sa0_s10));
  `include "b1.logic.vh"
endmodule

