// Test type: Hex Numbers - underscore within size
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=1_6'hC2d3;
endmodule
