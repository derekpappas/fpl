//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : ddr_bridge_ctrl.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module ddr_bridge_ctrl(dc_dbdummy5);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 27
  input dc_dbdummy5;
  `include "ddr_bridge_ctrl.logic.v"
endmodule

