// Test type: procedural continuous assignment - deassign variable lvalue
// Vparser rule name:
// Author: andreib
module procedural_continuous_assignment2;
reg a;
initial deassign a;
endmodule
