-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./b1_cslc_generated/code/vhdl/a1.vhd
-- FILE GENERATED ON : Wed Apr 29 21:51:03 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \a1\ is
  port(\p1\ : out csl_bit_vector(10#4# - 10#1# downto 10#0#));
begin
end entity;

architecture \a1_logic\ of \a1\ is
begin
end architecture;

