// Test type: Continuous assignment - h0, st1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous631;
wire a;
assign (highz0, strong1) a=1'b1;
endmodule
