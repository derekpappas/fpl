// Test type: always statement - nonblocking_assignment - no attribute instance
// Vparser rule name:
// Author: andreib
module alwcon19;
reg [7:0]a;
always a<=2;
endmodule
