module testbench_event_declaration;
    event_declaration0 event_declaration_instance0();
    event_declaration1 event_declaration_instance1();
    event_declaration2 event_declaration_instance2();
    event_declaration3 event_declaration_instance3();
    event_declaration4 event_declaration_instance4();
    event_declaration5 event_declaration_instance5();
    event_declaration6 event_declaration_instance6();
    event_declaration7 event_declaration_instance7();
    event_declaration8 event_declaration_instance8();
    event_declaration9 event_declaration_instance9();
    event_declaration10 event_declaration_instance10();
    event_declaration11 event_declaration_instance11();
    event_declaration12 event_declaration_instance12();
    event_declaration13 event_declaration_instance13();
    event_declaration14 event_declaration_instance14();
    event_declaration15 event_declaration_instance15();
    event_declaration16 event_declaration_instance16();
    event_declaration17 event_declaration_instance17();
    event_declaration18 event_declaration_instance18();
    event_declaration19 event_declaration_instance19();
    event_declaration20 event_declaration_instance20();
    event_declaration21 event_declaration_instance21();
    event_declaration22 event_declaration_instance22();
    event_declaration23 event_declaration_instance23();
    event_declaration24 event_declaration_instance24();
    event_declaration25 event_declaration_instance25();
    event_declaration26 event_declaration_instance26();
    event_declaration27 event_declaration_instance27();
    event_declaration28 event_declaration_instance28();
    event_declaration29 event_declaration_instance29();
    event_declaration30 event_declaration_instance30();
    event_declaration31 event_declaration_instance31();
    event_declaration32 event_declaration_instance32();
    event_declaration33 event_declaration_instance33();
    event_declaration34 event_declaration_instance34();
    event_declaration35 event_declaration_instance35();
    event_declaration36 event_declaration_instance36();
    event_declaration37 event_declaration_instance37();
    event_declaration38 event_declaration_instance38();
    event_declaration39 event_declaration_instance39();
    event_declaration40 event_declaration_instance40();
    event_declaration41 event_declaration_instance41();
    event_declaration42 event_declaration_instance42();
    event_declaration43 event_declaration_instance43();
    event_declaration44 event_declaration_instance44();
    event_declaration45 event_declaration_instance45();
    event_declaration46 event_declaration_instance46();
    event_declaration47 event_declaration_instance47();
    event_declaration48 event_declaration_instance48();
    event_declaration49 event_declaration_instance49();
    event_declaration50 event_declaration_instance50();
    event_declaration51 event_declaration_instance51();
    event_declaration52 event_declaration_instance52();
    event_declaration53 event_declaration_instance53();
    event_declaration54 event_declaration_instance54();
    event_declaration55 event_declaration_instance55();
    event_declaration56 event_declaration_instance56();
    event_declaration57 event_declaration_instance57();
    event_declaration58 event_declaration_instance58();
    event_declaration59 event_declaration_instance59();
    event_declaration60 event_declaration_instance60();
    event_declaration61 event_declaration_instance61();
    event_declaration62 event_declaration_instance62();
    event_declaration63 event_declaration_instance63();
    event_declaration64 event_declaration_instance64();
    event_declaration65 event_declaration_instance65();
    event_declaration66 event_declaration_instance66();
    event_declaration67 event_declaration_instance67();
    event_declaration68 event_declaration_instance68();
    event_declaration69 event_declaration_instance69();
    event_declaration70 event_declaration_instance70();
    event_declaration71 event_declaration_instance71();
    event_declaration72 event_declaration_instance72();
    event_declaration73 event_declaration_instance73();
    event_declaration74 event_declaration_instance74();
    event_declaration75 event_declaration_instance75();
    event_declaration76 event_declaration_instance76();
    event_declaration77 event_declaration_instance77();
    event_declaration78 event_declaration_instance78();
    event_declaration79 event_declaration_instance79();
    event_declaration80 event_declaration_instance80();
    event_declaration81 event_declaration_instance81();
    event_declaration82 event_declaration_instance82();
    event_declaration83 event_declaration_instance83();
endmodule
//@
//author : andreib
module event_declaration0;
event abc;
endmodule
//author : andreib
module event_declaration1;
event abc , ABC;
endmodule
//author : andreib
module event_declaration2;
event abc , ABC , _12;
endmodule
//author : andreib
module event_declaration3;
event abc , ABC , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration4;
event abc , ABC , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration5;
event abc , ABC , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration6;
event abc , ABC [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration7;
event abc , ABC [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration8;
event abc , ABC [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration9;
event abc , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration10;
event abc , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration11;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration12;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration13;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration14;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration15;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration16;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration17;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration18;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration19;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration20;
event abc , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration21;
event abc [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration22;
event abc [ 2 : 2 ] , ABC;
endmodule
//author : andreib
module event_declaration23;
event abc [ 2 : 2 ] , ABC , _12;
endmodule
//author : andreib
module event_declaration24;
event abc [ 2 : 2 ] , ABC , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration25;
event abc [ 2 : 2 ] , ABC , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration26;
event abc [ 2 : 2 ] , ABC , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration27;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration28;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration29;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration30;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration31;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration32;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration33;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration34;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration35;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration36;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration37;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration38;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration39;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration40;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration41;
event abc [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration42;
event abc [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration43;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC;
endmodule
//author : andreib
module event_declaration44;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC , _12;
endmodule
//author : andreib
module event_declaration45;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration46;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration47;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration48;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration49;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration50;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration51;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration52;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration53;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration54;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration55;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration56;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration57;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration58;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration59;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration60;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration61;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration62;
event abc [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration63;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration64;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC;
endmodule
//author : andreib
module event_declaration65;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC , _12;
endmodule
//author : andreib
module event_declaration66;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration67;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration68;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration69;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration70;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration71;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration72;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration73;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration74;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration75;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration76;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration77;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration78;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration79;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration80;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12;
endmodule
//author : andreib
module event_declaration81;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration82;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module event_declaration83;
event abc [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABC [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _12 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
