// Test type: Octal Numbers - no size lower case base
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a='O7460;
endmodule
