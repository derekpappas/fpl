// Test type: delay_control - delay_value - unsigned number
// Vparser rule name:
// Author: andreib
module delay_control1;
reg a;
initial #10 a=1'b1;
endmodule
