u4.vhd
