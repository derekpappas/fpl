// Test type: Binary Numbers - size and upper case base
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=3'B101;
endmodule
