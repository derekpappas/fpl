//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : dp_fp32_gasket.v
//FILE GENERATED ON : Tue Aug 12 09:34:23 2008

`include "defines.v"

module dp_fp32_gasket();
// Location of source csl unit: file name = generated/agent_cl.csl line number = 96
  `include "dp_fp32_gasket.logic.v"
endmodule

