`include "defines.v"

module s0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 127
  input [1 - 1:0] ar_sa0_s10;
  r0 r0(.ar_sa0_s10(ar_sa0_s10));
  `include "s0.logic.vh"
endmodule

