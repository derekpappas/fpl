// Test type: net_assignment - conditional expression
// Vparser rule name:
// Author: andreib
module netasign8;
wire a,b,c,d;
assign a=b?c:d;
endmodule
