module x;
   reg _389000_389000 ; 
   reg __389000_389000;
   reg _389001_389001 ; 
   reg __389001_389001;
   reg _389002_389002 ; 
   reg __389002_389002;
   reg _389003_389003 ; 
   reg __389003_389003;
   reg _389004_389004 ; 
   reg __389004_389004;
   reg _389005_389005 ; 
   reg __389005_389005;
   reg _389006_389006 ; 
   reg __389006_389006;
   reg _389007_389007 ; 
   reg __389007_389007;
   reg _389008_389008 ; 
   reg __389008_389008;
   reg _389009_389009 ; 
   reg __389009_389009;
   reg _389010_389010 ; 
   reg __389010_389010;
   reg _389011_389011 ; 
   reg __389011_389011;
   reg _389012_389012 ; 
   reg __389012_389012;
   reg _389013_389013 ; 
   reg __389013_389013;
   reg _389014_389014 ; 
   reg __389014_389014;
   reg _389015_389015 ; 
   reg __389015_389015;
   reg _389016_389016 ; 
   reg __389016_389016;
   reg _389017_389017 ; 
   reg __389017_389017;
   reg _389018_389018 ; 
   reg __389018_389018;
   reg _389019_389019 ; 
   reg __389019_389019;
   reg _389020_389020 ; 
   reg __389020_389020;
   reg _389021_389021 ; 
   reg __389021_389021;
   reg _389022_389022 ; 
   reg __389022_389022;
   reg _389023_389023 ; 
   reg __389023_389023;
   reg _389024_389024 ; 
   reg __389024_389024;
   reg _389025_389025 ; 
   reg __389025_389025;
   reg _389026_389026 ; 
   reg __389026_389026;
   reg _389027_389027 ; 
   reg __389027_389027;
   reg _389028_389028 ; 
   reg __389028_389028;
   reg _389029_389029 ; 
   reg __389029_389029;
   reg _389030_389030 ; 
   reg __389030_389030;
   reg _389031_389031 ; 
   reg __389031_389031;
   reg _389032_389032 ; 
   reg __389032_389032;
   reg _389033_389033 ; 
   reg __389033_389033;
   reg _389034_389034 ; 
   reg __389034_389034;
   reg _389035_389035 ; 
   reg __389035_389035;
   reg _389036_389036 ; 
   reg __389036_389036;
   reg _389037_389037 ; 
   reg __389037_389037;
   reg _389038_389038 ; 
   reg __389038_389038;
   reg _389039_389039 ; 
   reg __389039_389039;
   reg _389040_389040 ; 
   reg __389040_389040;
   reg _389041_389041 ; 
   reg __389041_389041;
   reg _389042_389042 ; 
   reg __389042_389042;
   reg _389043_389043 ; 
   reg __389043_389043;
   reg _389044_389044 ; 
   reg __389044_389044;
   reg _389045_389045 ; 
   reg __389045_389045;
   reg _389046_389046 ; 
   reg __389046_389046;
   reg _389047_389047 ; 
   reg __389047_389047;
   reg _389048_389048 ; 
   reg __389048_389048;
   reg _389049_389049 ; 
   reg __389049_389049;
   reg _389050_389050 ; 
   reg __389050_389050;
   reg _389051_389051 ; 
   reg __389051_389051;
   reg _389052_389052 ; 
   reg __389052_389052;
   reg _389053_389053 ; 
   reg __389053_389053;
   reg _389054_389054 ; 
   reg __389054_389054;
   reg _389055_389055 ; 
   reg __389055_389055;
   reg _389056_389056 ; 
   reg __389056_389056;
   reg _389057_389057 ; 
   reg __389057_389057;
   reg _389058_389058 ; 
   reg __389058_389058;
   reg _389059_389059 ; 
   reg __389059_389059;
   reg _389060_389060 ; 
   reg __389060_389060;
   reg _389061_389061 ; 
   reg __389061_389061;
   reg _389062_389062 ; 
   reg __389062_389062;
   reg _389063_389063 ; 
   reg __389063_389063;
   reg _389064_389064 ; 
   reg __389064_389064;
   reg _389065_389065 ; 
   reg __389065_389065;
   reg _389066_389066 ; 
   reg __389066_389066;
   reg _389067_389067 ; 
   reg __389067_389067;
   reg _389068_389068 ; 
   reg __389068_389068;
   reg _389069_389069 ; 
   reg __389069_389069;
   reg _389070_389070 ; 
   reg __389070_389070;
   reg _389071_389071 ; 
   reg __389071_389071;
   reg _389072_389072 ; 
   reg __389072_389072;
   reg _389073_389073 ; 
   reg __389073_389073;
   reg _389074_389074 ; 
   reg __389074_389074;
   reg _389075_389075 ; 
   reg __389075_389075;
   reg _389076_389076 ; 
   reg __389076_389076;
   reg _389077_389077 ; 
   reg __389077_389077;
   reg _389078_389078 ; 
   reg __389078_389078;
   reg _389079_389079 ; 
   reg __389079_389079;
   reg _389080_389080 ; 
   reg __389080_389080;
   reg _389081_389081 ; 
   reg __389081_389081;
   reg _389082_389082 ; 
   reg __389082_389082;
   reg _389083_389083 ; 
   reg __389083_389083;
   reg _389084_389084 ; 
   reg __389084_389084;
   reg _389085_389085 ; 
   reg __389085_389085;
   reg _389086_389086 ; 
   reg __389086_389086;
   reg _389087_389087 ; 
   reg __389087_389087;
   reg _389088_389088 ; 
   reg __389088_389088;
   reg _389089_389089 ; 
   reg __389089_389089;
   reg _389090_389090 ; 
   reg __389090_389090;
   reg _389091_389091 ; 
   reg __389091_389091;
   reg _389092_389092 ; 
   reg __389092_389092;
   reg _389093_389093 ; 
   reg __389093_389093;
   reg _389094_389094 ; 
   reg __389094_389094;
   reg _389095_389095 ; 
   reg __389095_389095;
   reg _389096_389096 ; 
   reg __389096_389096;
   reg _389097_389097 ; 
   reg __389097_389097;
   reg _389098_389098 ; 
   reg __389098_389098;
   reg _389099_389099 ; 
   reg __389099_389099;
   reg _389100_389100 ; 
   reg __389100_389100;
   reg _389101_389101 ; 
   reg __389101_389101;
   reg _389102_389102 ; 
   reg __389102_389102;
   reg _389103_389103 ; 
   reg __389103_389103;
   reg _389104_389104 ; 
   reg __389104_389104;
   reg _389105_389105 ; 
   reg __389105_389105;
   reg _389106_389106 ; 
   reg __389106_389106;
   reg _389107_389107 ; 
   reg __389107_389107;
   reg _389108_389108 ; 
   reg __389108_389108;
   reg _389109_389109 ; 
   reg __389109_389109;
   reg _389110_389110 ; 
   reg __389110_389110;
   reg _389111_389111 ; 
   reg __389111_389111;
   reg _389112_389112 ; 
   reg __389112_389112;
   reg _389113_389113 ; 
   reg __389113_389113;
   reg _389114_389114 ; 
   reg __389114_389114;
   reg _389115_389115 ; 
   reg __389115_389115;
   reg _389116_389116 ; 
   reg __389116_389116;
   reg _389117_389117 ; 
   reg __389117_389117;
   reg _389118_389118 ; 
   reg __389118_389118;
   reg _389119_389119 ; 
   reg __389119_389119;
   reg _389120_389120 ; 
   reg __389120_389120;
   reg _389121_389121 ; 
   reg __389121_389121;
   reg _389122_389122 ; 
   reg __389122_389122;
   reg _389123_389123 ; 
   reg __389123_389123;
   reg _389124_389124 ; 
   reg __389124_389124;
   reg _389125_389125 ; 
   reg __389125_389125;
   reg _389126_389126 ; 
   reg __389126_389126;
   reg _389127_389127 ; 
   reg __389127_389127;
   reg _389128_389128 ; 
   reg __389128_389128;
   reg _389129_389129 ; 
   reg __389129_389129;
   reg _389130_389130 ; 
   reg __389130_389130;
   reg _389131_389131 ; 
   reg __389131_389131;
   reg _389132_389132 ; 
   reg __389132_389132;
   reg _389133_389133 ; 
   reg __389133_389133;
   reg _389134_389134 ; 
   reg __389134_389134;
   reg _389135_389135 ; 
   reg __389135_389135;
   reg _389136_389136 ; 
   reg __389136_389136;
   reg _389137_389137 ; 
   reg __389137_389137;
   reg _389138_389138 ; 
   reg __389138_389138;
   reg _389139_389139 ; 
   reg __389139_389139;
   reg _389140_389140 ; 
   reg __389140_389140;
   reg _389141_389141 ; 
   reg __389141_389141;
   reg _389142_389142 ; 
   reg __389142_389142;
   reg _389143_389143 ; 
   reg __389143_389143;
   reg _389144_389144 ; 
   reg __389144_389144;
   reg _389145_389145 ; 
   reg __389145_389145;
   reg _389146_389146 ; 
   reg __389146_389146;
   reg _389147_389147 ; 
   reg __389147_389147;
   reg _389148_389148 ; 
   reg __389148_389148;
   reg _389149_389149 ; 
   reg __389149_389149;
   reg _389150_389150 ; 
   reg __389150_389150;
   reg _389151_389151 ; 
   reg __389151_389151;
   reg _389152_389152 ; 
   reg __389152_389152;
   reg _389153_389153 ; 
   reg __389153_389153;
   reg _389154_389154 ; 
   reg __389154_389154;
   reg _389155_389155 ; 
   reg __389155_389155;
   reg _389156_389156 ; 
   reg __389156_389156;
   reg _389157_389157 ; 
   reg __389157_389157;
   reg _389158_389158 ; 
   reg __389158_389158;
   reg _389159_389159 ; 
   reg __389159_389159;
   reg _389160_389160 ; 
   reg __389160_389160;
   reg _389161_389161 ; 
   reg __389161_389161;
   reg _389162_389162 ; 
   reg __389162_389162;
   reg _389163_389163 ; 
   reg __389163_389163;
   reg _389164_389164 ; 
   reg __389164_389164;
   reg _389165_389165 ; 
   reg __389165_389165;
   reg _389166_389166 ; 
   reg __389166_389166;
   reg _389167_389167 ; 
   reg __389167_389167;
   reg _389168_389168 ; 
   reg __389168_389168;
   reg _389169_389169 ; 
   reg __389169_389169;
   reg _389170_389170 ; 
   reg __389170_389170;
   reg _389171_389171 ; 
   reg __389171_389171;
   reg _389172_389172 ; 
   reg __389172_389172;
   reg _389173_389173 ; 
   reg __389173_389173;
   reg _389174_389174 ; 
   reg __389174_389174;
   reg _389175_389175 ; 
   reg __389175_389175;
   reg _389176_389176 ; 
   reg __389176_389176;
   reg _389177_389177 ; 
   reg __389177_389177;
   reg _389178_389178 ; 
   reg __389178_389178;
   reg _389179_389179 ; 
   reg __389179_389179;
   reg _389180_389180 ; 
   reg __389180_389180;
   reg _389181_389181 ; 
   reg __389181_389181;
   reg _389182_389182 ; 
   reg __389182_389182;
   reg _389183_389183 ; 
   reg __389183_389183;
   reg _389184_389184 ; 
   reg __389184_389184;
   reg _389185_389185 ; 
   reg __389185_389185;
   reg _389186_389186 ; 
   reg __389186_389186;
   reg _389187_389187 ; 
   reg __389187_389187;
   reg _389188_389188 ; 
   reg __389188_389188;
   reg _389189_389189 ; 
   reg __389189_389189;
   reg _389190_389190 ; 
   reg __389190_389190;
   reg _389191_389191 ; 
   reg __389191_389191;
   reg _389192_389192 ; 
   reg __389192_389192;
   reg _389193_389193 ; 
   reg __389193_389193;
   reg _389194_389194 ; 
   reg __389194_389194;
   reg _389195_389195 ; 
   reg __389195_389195;
   reg _389196_389196 ; 
   reg __389196_389196;
   reg _389197_389197 ; 
   reg __389197_389197;
   reg _389198_389198 ; 
   reg __389198_389198;
   reg _389199_389199 ; 
   reg __389199_389199;
   reg _389200_389200 ; 
   reg __389200_389200;
   reg _389201_389201 ; 
   reg __389201_389201;
   reg _389202_389202 ; 
   reg __389202_389202;
   reg _389203_389203 ; 
   reg __389203_389203;
   reg _389204_389204 ; 
   reg __389204_389204;
   reg _389205_389205 ; 
   reg __389205_389205;
   reg _389206_389206 ; 
   reg __389206_389206;
   reg _389207_389207 ; 
   reg __389207_389207;
   reg _389208_389208 ; 
   reg __389208_389208;
   reg _389209_389209 ; 
   reg __389209_389209;
   reg _389210_389210 ; 
   reg __389210_389210;
   reg _389211_389211 ; 
   reg __389211_389211;
   reg _389212_389212 ; 
   reg __389212_389212;
   reg _389213_389213 ; 
   reg __389213_389213;
   reg _389214_389214 ; 
   reg __389214_389214;
   reg _389215_389215 ; 
   reg __389215_389215;
   reg _389216_389216 ; 
   reg __389216_389216;
   reg _389217_389217 ; 
   reg __389217_389217;
   reg _389218_389218 ; 
   reg __389218_389218;
   reg _389219_389219 ; 
   reg __389219_389219;
   reg _389220_389220 ; 
   reg __389220_389220;
   reg _389221_389221 ; 
   reg __389221_389221;
   reg _389222_389222 ; 
   reg __389222_389222;
   reg _389223_389223 ; 
   reg __389223_389223;
   reg _389224_389224 ; 
   reg __389224_389224;
   reg _389225_389225 ; 
   reg __389225_389225;
   reg _389226_389226 ; 
   reg __389226_389226;
   reg _389227_389227 ; 
   reg __389227_389227;
   reg _389228_389228 ; 
   reg __389228_389228;
   reg _389229_389229 ; 
   reg __389229_389229;
   reg _389230_389230 ; 
   reg __389230_389230;
   reg _389231_389231 ; 
   reg __389231_389231;
   reg _389232_389232 ; 
   reg __389232_389232;
   reg _389233_389233 ; 
   reg __389233_389233;
   reg _389234_389234 ; 
   reg __389234_389234;
   reg _389235_389235 ; 
   reg __389235_389235;
   reg _389236_389236 ; 
   reg __389236_389236;
   reg _389237_389237 ; 
   reg __389237_389237;
   reg _389238_389238 ; 
   reg __389238_389238;
   reg _389239_389239 ; 
   reg __389239_389239;
   reg _389240_389240 ; 
   reg __389240_389240;
   reg _389241_389241 ; 
   reg __389241_389241;
   reg _389242_389242 ; 
   reg __389242_389242;
   reg _389243_389243 ; 
   reg __389243_389243;
   reg _389244_389244 ; 
   reg __389244_389244;
   reg _389245_389245 ; 
   reg __389245_389245;
   reg _389246_389246 ; 
   reg __389246_389246;
   reg _389247_389247 ; 
   reg __389247_389247;
   reg _389248_389248 ; 
   reg __389248_389248;
   reg _389249_389249 ; 
   reg __389249_389249;
   reg _389250_389250 ; 
   reg __389250_389250;
   reg _389251_389251 ; 
   reg __389251_389251;
   reg _389252_389252 ; 
   reg __389252_389252;
   reg _389253_389253 ; 
   reg __389253_389253;
   reg _389254_389254 ; 
   reg __389254_389254;
   reg _389255_389255 ; 
   reg __389255_389255;
   reg _389256_389256 ; 
   reg __389256_389256;
   reg _389257_389257 ; 
   reg __389257_389257;
   reg _389258_389258 ; 
   reg __389258_389258;
   reg _389259_389259 ; 
   reg __389259_389259;
   reg _389260_389260 ; 
   reg __389260_389260;
   reg _389261_389261 ; 
   reg __389261_389261;
   reg _389262_389262 ; 
   reg __389262_389262;
   reg _389263_389263 ; 
   reg __389263_389263;
   reg _389264_389264 ; 
   reg __389264_389264;
   reg _389265_389265 ; 
   reg __389265_389265;
   reg _389266_389266 ; 
   reg __389266_389266;
   reg _389267_389267 ; 
   reg __389267_389267;
   reg _389268_389268 ; 
   reg __389268_389268;
   reg _389269_389269 ; 
   reg __389269_389269;
   reg _389270_389270 ; 
   reg __389270_389270;
   reg _389271_389271 ; 
   reg __389271_389271;
   reg _389272_389272 ; 
   reg __389272_389272;
   reg _389273_389273 ; 
   reg __389273_389273;
   reg _389274_389274 ; 
   reg __389274_389274;
   reg _389275_389275 ; 
   reg __389275_389275;
   reg _389276_389276 ; 
   reg __389276_389276;
   reg _389277_389277 ; 
   reg __389277_389277;
   reg _389278_389278 ; 
   reg __389278_389278;
   reg _389279_389279 ; 
   reg __389279_389279;
   reg _389280_389280 ; 
   reg __389280_389280;
   reg _389281_389281 ; 
   reg __389281_389281;
   reg _389282_389282 ; 
   reg __389282_389282;
   reg _389283_389283 ; 
   reg __389283_389283;
   reg _389284_389284 ; 
   reg __389284_389284;
   reg _389285_389285 ; 
   reg __389285_389285;
   reg _389286_389286 ; 
   reg __389286_389286;
   reg _389287_389287 ; 
   reg __389287_389287;
   reg _389288_389288 ; 
   reg __389288_389288;
   reg _389289_389289 ; 
   reg __389289_389289;
   reg _389290_389290 ; 
   reg __389290_389290;
   reg _389291_389291 ; 
   reg __389291_389291;
   reg _389292_389292 ; 
   reg __389292_389292;
   reg _389293_389293 ; 
   reg __389293_389293;
   reg _389294_389294 ; 
   reg __389294_389294;
   reg _389295_389295 ; 
   reg __389295_389295;
   reg _389296_389296 ; 
   reg __389296_389296;
   reg _389297_389297 ; 
   reg __389297_389297;
   reg _389298_389298 ; 
   reg __389298_389298;
   reg _389299_389299 ; 
   reg __389299_389299;
   reg _389300_389300 ; 
   reg __389300_389300;
   reg _389301_389301 ; 
   reg __389301_389301;
   reg _389302_389302 ; 
   reg __389302_389302;
   reg _389303_389303 ; 
   reg __389303_389303;
   reg _389304_389304 ; 
   reg __389304_389304;
   reg _389305_389305 ; 
   reg __389305_389305;
   reg _389306_389306 ; 
   reg __389306_389306;
   reg _389307_389307 ; 
   reg __389307_389307;
   reg _389308_389308 ; 
   reg __389308_389308;
   reg _389309_389309 ; 
   reg __389309_389309;
   reg _389310_389310 ; 
   reg __389310_389310;
   reg _389311_389311 ; 
   reg __389311_389311;
   reg _389312_389312 ; 
   reg __389312_389312;
   reg _389313_389313 ; 
   reg __389313_389313;
   reg _389314_389314 ; 
   reg __389314_389314;
   reg _389315_389315 ; 
   reg __389315_389315;
   reg _389316_389316 ; 
   reg __389316_389316;
   reg _389317_389317 ; 
   reg __389317_389317;
   reg _389318_389318 ; 
   reg __389318_389318;
   reg _389319_389319 ; 
   reg __389319_389319;
   reg _389320_389320 ; 
   reg __389320_389320;
   reg _389321_389321 ; 
   reg __389321_389321;
   reg _389322_389322 ; 
   reg __389322_389322;
   reg _389323_389323 ; 
   reg __389323_389323;
   reg _389324_389324 ; 
   reg __389324_389324;
   reg _389325_389325 ; 
   reg __389325_389325;
   reg _389326_389326 ; 
   reg __389326_389326;
   reg _389327_389327 ; 
   reg __389327_389327;
   reg _389328_389328 ; 
   reg __389328_389328;
   reg _389329_389329 ; 
   reg __389329_389329;
   reg _389330_389330 ; 
   reg __389330_389330;
   reg _389331_389331 ; 
   reg __389331_389331;
   reg _389332_389332 ; 
   reg __389332_389332;
   reg _389333_389333 ; 
   reg __389333_389333;
   reg _389334_389334 ; 
   reg __389334_389334;
   reg _389335_389335 ; 
   reg __389335_389335;
   reg _389336_389336 ; 
   reg __389336_389336;
   reg _389337_389337 ; 
   reg __389337_389337;
   reg _389338_389338 ; 
   reg __389338_389338;
   reg _389339_389339 ; 
   reg __389339_389339;
   reg _389340_389340 ; 
   reg __389340_389340;
   reg _389341_389341 ; 
   reg __389341_389341;
   reg _389342_389342 ; 
   reg __389342_389342;
   reg _389343_389343 ; 
   reg __389343_389343;
   reg _389344_389344 ; 
   reg __389344_389344;
   reg _389345_389345 ; 
   reg __389345_389345;
   reg _389346_389346 ; 
   reg __389346_389346;
   reg _389347_389347 ; 
   reg __389347_389347;
   reg _389348_389348 ; 
   reg __389348_389348;
   reg _389349_389349 ; 
   reg __389349_389349;
   reg _389350_389350 ; 
   reg __389350_389350;
   reg _389351_389351 ; 
   reg __389351_389351;
   reg _389352_389352 ; 
   reg __389352_389352;
   reg _389353_389353 ; 
   reg __389353_389353;
   reg _389354_389354 ; 
   reg __389354_389354;
   reg _389355_389355 ; 
   reg __389355_389355;
   reg _389356_389356 ; 
   reg __389356_389356;
   reg _389357_389357 ; 
   reg __389357_389357;
   reg _389358_389358 ; 
   reg __389358_389358;
   reg _389359_389359 ; 
   reg __389359_389359;
   reg _389360_389360 ; 
   reg __389360_389360;
   reg _389361_389361 ; 
   reg __389361_389361;
   reg _389362_389362 ; 
   reg __389362_389362;
   reg _389363_389363 ; 
   reg __389363_389363;
   reg _389364_389364 ; 
   reg __389364_389364;
   reg _389365_389365 ; 
   reg __389365_389365;
   reg _389366_389366 ; 
   reg __389366_389366;
   reg _389367_389367 ; 
   reg __389367_389367;
   reg _389368_389368 ; 
   reg __389368_389368;
   reg _389369_389369 ; 
   reg __389369_389369;
   reg _389370_389370 ; 
   reg __389370_389370;
   reg _389371_389371 ; 
   reg __389371_389371;
   reg _389372_389372 ; 
   reg __389372_389372;
   reg _389373_389373 ; 
   reg __389373_389373;
   reg _389374_389374 ; 
   reg __389374_389374;
   reg _389375_389375 ; 
   reg __389375_389375;
   reg _389376_389376 ; 
   reg __389376_389376;
   reg _389377_389377 ; 
   reg __389377_389377;
   reg _389378_389378 ; 
   reg __389378_389378;
   reg _389379_389379 ; 
   reg __389379_389379;
   reg _389380_389380 ; 
   reg __389380_389380;
   reg _389381_389381 ; 
   reg __389381_389381;
   reg _389382_389382 ; 
   reg __389382_389382;
   reg _389383_389383 ; 
   reg __389383_389383;
   reg _389384_389384 ; 
   reg __389384_389384;
   reg _389385_389385 ; 
   reg __389385_389385;
   reg _389386_389386 ; 
   reg __389386_389386;
   reg _389387_389387 ; 
   reg __389387_389387;
   reg _389388_389388 ; 
   reg __389388_389388;
   reg _389389_389389 ; 
   reg __389389_389389;
   reg _389390_389390 ; 
   reg __389390_389390;
   reg _389391_389391 ; 
   reg __389391_389391;
   reg _389392_389392 ; 
   reg __389392_389392;
   reg _389393_389393 ; 
   reg __389393_389393;
   reg _389394_389394 ; 
   reg __389394_389394;
   reg _389395_389395 ; 
   reg __389395_389395;
   reg _389396_389396 ; 
   reg __389396_389396;
   reg _389397_389397 ; 
   reg __389397_389397;
   reg _389398_389398 ; 
   reg __389398_389398;
   reg _389399_389399 ; 
   reg __389399_389399;
   reg _389400_389400 ; 
   reg __389400_389400;
   reg _389401_389401 ; 
   reg __389401_389401;
   reg _389402_389402 ; 
   reg __389402_389402;
   reg _389403_389403 ; 
   reg __389403_389403;
   reg _389404_389404 ; 
   reg __389404_389404;
   reg _389405_389405 ; 
   reg __389405_389405;
   reg _389406_389406 ; 
   reg __389406_389406;
   reg _389407_389407 ; 
   reg __389407_389407;
   reg _389408_389408 ; 
   reg __389408_389408;
   reg _389409_389409 ; 
   reg __389409_389409;
   reg _389410_389410 ; 
   reg __389410_389410;
   reg _389411_389411 ; 
   reg __389411_389411;
   reg _389412_389412 ; 
   reg __389412_389412;
   reg _389413_389413 ; 
   reg __389413_389413;
   reg _389414_389414 ; 
   reg __389414_389414;
   reg _389415_389415 ; 
   reg __389415_389415;
   reg _389416_389416 ; 
   reg __389416_389416;
   reg _389417_389417 ; 
   reg __389417_389417;
   reg _389418_389418 ; 
   reg __389418_389418;
   reg _389419_389419 ; 
   reg __389419_389419;
   reg _389420_389420 ; 
   reg __389420_389420;
   reg _389421_389421 ; 
   reg __389421_389421;
   reg _389422_389422 ; 
   reg __389422_389422;
   reg _389423_389423 ; 
   reg __389423_389423;
   reg _389424_389424 ; 
   reg __389424_389424;
   reg _389425_389425 ; 
   reg __389425_389425;
   reg _389426_389426 ; 
   reg __389426_389426;
   reg _389427_389427 ; 
   reg __389427_389427;
   reg _389428_389428 ; 
   reg __389428_389428;
   reg _389429_389429 ; 
   reg __389429_389429;
   reg _389430_389430 ; 
   reg __389430_389430;
   reg _389431_389431 ; 
   reg __389431_389431;
   reg _389432_389432 ; 
   reg __389432_389432;
   reg _389433_389433 ; 
   reg __389433_389433;
   reg _389434_389434 ; 
   reg __389434_389434;
   reg _389435_389435 ; 
   reg __389435_389435;
   reg _389436_389436 ; 
   reg __389436_389436;
   reg _389437_389437 ; 
   reg __389437_389437;
   reg _389438_389438 ; 
   reg __389438_389438;
   reg _389439_389439 ; 
   reg __389439_389439;
   reg _389440_389440 ; 
   reg __389440_389440;
   reg _389441_389441 ; 
   reg __389441_389441;
   reg _389442_389442 ; 
   reg __389442_389442;
   reg _389443_389443 ; 
   reg __389443_389443;
   reg _389444_389444 ; 
   reg __389444_389444;
   reg _389445_389445 ; 
   reg __389445_389445;
   reg _389446_389446 ; 
   reg __389446_389446;
   reg _389447_389447 ; 
   reg __389447_389447;
   reg _389448_389448 ; 
   reg __389448_389448;
   reg _389449_389449 ; 
   reg __389449_389449;
   reg _389450_389450 ; 
   reg __389450_389450;
   reg _389451_389451 ; 
   reg __389451_389451;
   reg _389452_389452 ; 
   reg __389452_389452;
   reg _389453_389453 ; 
   reg __389453_389453;
   reg _389454_389454 ; 
   reg __389454_389454;
   reg _389455_389455 ; 
   reg __389455_389455;
   reg _389456_389456 ; 
   reg __389456_389456;
   reg _389457_389457 ; 
   reg __389457_389457;
   reg _389458_389458 ; 
   reg __389458_389458;
   reg _389459_389459 ; 
   reg __389459_389459;
   reg _389460_389460 ; 
   reg __389460_389460;
   reg _389461_389461 ; 
   reg __389461_389461;
   reg _389462_389462 ; 
   reg __389462_389462;
   reg _389463_389463 ; 
   reg __389463_389463;
   reg _389464_389464 ; 
   reg __389464_389464;
   reg _389465_389465 ; 
   reg __389465_389465;
   reg _389466_389466 ; 
   reg __389466_389466;
   reg _389467_389467 ; 
   reg __389467_389467;
   reg _389468_389468 ; 
   reg __389468_389468;
   reg _389469_389469 ; 
   reg __389469_389469;
   reg _389470_389470 ; 
   reg __389470_389470;
   reg _389471_389471 ; 
   reg __389471_389471;
   reg _389472_389472 ; 
   reg __389472_389472;
   reg _389473_389473 ; 
   reg __389473_389473;
   reg _389474_389474 ; 
   reg __389474_389474;
   reg _389475_389475 ; 
   reg __389475_389475;
   reg _389476_389476 ; 
   reg __389476_389476;
   reg _389477_389477 ; 
   reg __389477_389477;
   reg _389478_389478 ; 
   reg __389478_389478;
   reg _389479_389479 ; 
   reg __389479_389479;
   reg _389480_389480 ; 
   reg __389480_389480;
   reg _389481_389481 ; 
   reg __389481_389481;
   reg _389482_389482 ; 
   reg __389482_389482;
   reg _389483_389483 ; 
   reg __389483_389483;
   reg _389484_389484 ; 
   reg __389484_389484;
   reg _389485_389485 ; 
   reg __389485_389485;
   reg _389486_389486 ; 
   reg __389486_389486;
   reg _389487_389487 ; 
   reg __389487_389487;
   reg _389488_389488 ; 
   reg __389488_389488;
   reg _389489_389489 ; 
   reg __389489_389489;
   reg _389490_389490 ; 
   reg __389490_389490;
   reg _389491_389491 ; 
   reg __389491_389491;
   reg _389492_389492 ; 
   reg __389492_389492;
   reg _389493_389493 ; 
   reg __389493_389493;
   reg _389494_389494 ; 
   reg __389494_389494;
   reg _389495_389495 ; 
   reg __389495_389495;
   reg _389496_389496 ; 
   reg __389496_389496;
   reg _389497_389497 ; 
   reg __389497_389497;
   reg _389498_389498 ; 
   reg __389498_389498;
   reg _389499_389499 ; 
   reg __389499_389499;
   reg _389500_389500 ; 
   reg __389500_389500;
   reg _389501_389501 ; 
   reg __389501_389501;
   reg _389502_389502 ; 
   reg __389502_389502;
   reg _389503_389503 ; 
   reg __389503_389503;
   reg _389504_389504 ; 
   reg __389504_389504;
   reg _389505_389505 ; 
   reg __389505_389505;
   reg _389506_389506 ; 
   reg __389506_389506;
   reg _389507_389507 ; 
   reg __389507_389507;
   reg _389508_389508 ; 
   reg __389508_389508;
   reg _389509_389509 ; 
   reg __389509_389509;
   reg _389510_389510 ; 
   reg __389510_389510;
   reg _389511_389511 ; 
   reg __389511_389511;
   reg _389512_389512 ; 
   reg __389512_389512;
   reg _389513_389513 ; 
   reg __389513_389513;
   reg _389514_389514 ; 
   reg __389514_389514;
   reg _389515_389515 ; 
   reg __389515_389515;
   reg _389516_389516 ; 
   reg __389516_389516;
   reg _389517_389517 ; 
   reg __389517_389517;
   reg _389518_389518 ; 
   reg __389518_389518;
   reg _389519_389519 ; 
   reg __389519_389519;
   reg _389520_389520 ; 
   reg __389520_389520;
   reg _389521_389521 ; 
   reg __389521_389521;
   reg _389522_389522 ; 
   reg __389522_389522;
   reg _389523_389523 ; 
   reg __389523_389523;
   reg _389524_389524 ; 
   reg __389524_389524;
   reg _389525_389525 ; 
   reg __389525_389525;
   reg _389526_389526 ; 
   reg __389526_389526;
   reg _389527_389527 ; 
   reg __389527_389527;
   reg _389528_389528 ; 
   reg __389528_389528;
   reg _389529_389529 ; 
   reg __389529_389529;
   reg _389530_389530 ; 
   reg __389530_389530;
   reg _389531_389531 ; 
   reg __389531_389531;
   reg _389532_389532 ; 
   reg __389532_389532;
   reg _389533_389533 ; 
   reg __389533_389533;
   reg _389534_389534 ; 
   reg __389534_389534;
   reg _389535_389535 ; 
   reg __389535_389535;
   reg _389536_389536 ; 
   reg __389536_389536;
   reg _389537_389537 ; 
   reg __389537_389537;
   reg _389538_389538 ; 
   reg __389538_389538;
   reg _389539_389539 ; 
   reg __389539_389539;
   reg _389540_389540 ; 
   reg __389540_389540;
   reg _389541_389541 ; 
   reg __389541_389541;
   reg _389542_389542 ; 
   reg __389542_389542;
   reg _389543_389543 ; 
   reg __389543_389543;
   reg _389544_389544 ; 
   reg __389544_389544;
   reg _389545_389545 ; 
   reg __389545_389545;
   reg _389546_389546 ; 
   reg __389546_389546;
   reg _389547_389547 ; 
   reg __389547_389547;
   reg _389548_389548 ; 
   reg __389548_389548;
   reg _389549_389549 ; 
   reg __389549_389549;
   reg _389550_389550 ; 
   reg __389550_389550;
   reg _389551_389551 ; 
   reg __389551_389551;
   reg _389552_389552 ; 
   reg __389552_389552;
   reg _389553_389553 ; 
   reg __389553_389553;
   reg _389554_389554 ; 
   reg __389554_389554;
   reg _389555_389555 ; 
   reg __389555_389555;
   reg _389556_389556 ; 
   reg __389556_389556;
   reg _389557_389557 ; 
   reg __389557_389557;
   reg _389558_389558 ; 
   reg __389558_389558;
   reg _389559_389559 ; 
   reg __389559_389559;
   reg _389560_389560 ; 
   reg __389560_389560;
   reg _389561_389561 ; 
   reg __389561_389561;
   reg _389562_389562 ; 
   reg __389562_389562;
   reg _389563_389563 ; 
   reg __389563_389563;
   reg _389564_389564 ; 
   reg __389564_389564;
   reg _389565_389565 ; 
   reg __389565_389565;
   reg _389566_389566 ; 
   reg __389566_389566;
   reg _389567_389567 ; 
   reg __389567_389567;
   reg _389568_389568 ; 
   reg __389568_389568;
   reg _389569_389569 ; 
   reg __389569_389569;
   reg _389570_389570 ; 
   reg __389570_389570;
   reg _389571_389571 ; 
   reg __389571_389571;
   reg _389572_389572 ; 
   reg __389572_389572;
   reg _389573_389573 ; 
   reg __389573_389573;
   reg _389574_389574 ; 
   reg __389574_389574;
   reg _389575_389575 ; 
   reg __389575_389575;
   reg _389576_389576 ; 
   reg __389576_389576;
   reg _389577_389577 ; 
   reg __389577_389577;
   reg _389578_389578 ; 
   reg __389578_389578;
   reg _389579_389579 ; 
   reg __389579_389579;
   reg _389580_389580 ; 
   reg __389580_389580;
   reg _389581_389581 ; 
   reg __389581_389581;
   reg _389582_389582 ; 
   reg __389582_389582;
   reg _389583_389583 ; 
   reg __389583_389583;
   reg _389584_389584 ; 
   reg __389584_389584;
   reg _389585_389585 ; 
   reg __389585_389585;
   reg _389586_389586 ; 
   reg __389586_389586;
   reg _389587_389587 ; 
   reg __389587_389587;
   reg _389588_389588 ; 
   reg __389588_389588;
   reg _389589_389589 ; 
   reg __389589_389589;
   reg _389590_389590 ; 
   reg __389590_389590;
   reg _389591_389591 ; 
   reg __389591_389591;
   reg _389592_389592 ; 
   reg __389592_389592;
   reg _389593_389593 ; 
   reg __389593_389593;
   reg _389594_389594 ; 
   reg __389594_389594;
   reg _389595_389595 ; 
   reg __389595_389595;
   reg _389596_389596 ; 
   reg __389596_389596;
   reg _389597_389597 ; 
   reg __389597_389597;
   reg _389598_389598 ; 
   reg __389598_389598;
   reg _389599_389599 ; 
   reg __389599_389599;
   reg _389600_389600 ; 
   reg __389600_389600;
   reg _389601_389601 ; 
   reg __389601_389601;
   reg _389602_389602 ; 
   reg __389602_389602;
   reg _389603_389603 ; 
   reg __389603_389603;
   reg _389604_389604 ; 
   reg __389604_389604;
   reg _389605_389605 ; 
   reg __389605_389605;
   reg _389606_389606 ; 
   reg __389606_389606;
   reg _389607_389607 ; 
   reg __389607_389607;
   reg _389608_389608 ; 
   reg __389608_389608;
   reg _389609_389609 ; 
   reg __389609_389609;
   reg _389610_389610 ; 
   reg __389610_389610;
   reg _389611_389611 ; 
   reg __389611_389611;
   reg _389612_389612 ; 
   reg __389612_389612;
   reg _389613_389613 ; 
   reg __389613_389613;
   reg _389614_389614 ; 
   reg __389614_389614;
   reg _389615_389615 ; 
   reg __389615_389615;
   reg _389616_389616 ; 
   reg __389616_389616;
   reg _389617_389617 ; 
   reg __389617_389617;
   reg _389618_389618 ; 
   reg __389618_389618;
   reg _389619_389619 ; 
   reg __389619_389619;
   reg _389620_389620 ; 
   reg __389620_389620;
   reg _389621_389621 ; 
   reg __389621_389621;
   reg _389622_389622 ; 
   reg __389622_389622;
   reg _389623_389623 ; 
   reg __389623_389623;
   reg _389624_389624 ; 
   reg __389624_389624;
   reg _389625_389625 ; 
   reg __389625_389625;
   reg _389626_389626 ; 
   reg __389626_389626;
   reg _389627_389627 ; 
   reg __389627_389627;
   reg _389628_389628 ; 
   reg __389628_389628;
   reg _389629_389629 ; 
   reg __389629_389629;
   reg _389630_389630 ; 
   reg __389630_389630;
   reg _389631_389631 ; 
   reg __389631_389631;
   reg _389632_389632 ; 
   reg __389632_389632;
   reg _389633_389633 ; 
   reg __389633_389633;
   reg _389634_389634 ; 
   reg __389634_389634;
   reg _389635_389635 ; 
   reg __389635_389635;
   reg _389636_389636 ; 
   reg __389636_389636;
   reg _389637_389637 ; 
   reg __389637_389637;
   reg _389638_389638 ; 
   reg __389638_389638;
   reg _389639_389639 ; 
   reg __389639_389639;
   reg _389640_389640 ; 
   reg __389640_389640;
   reg _389641_389641 ; 
   reg __389641_389641;
   reg _389642_389642 ; 
   reg __389642_389642;
   reg _389643_389643 ; 
   reg __389643_389643;
   reg _389644_389644 ; 
   reg __389644_389644;
   reg _389645_389645 ; 
   reg __389645_389645;
   reg _389646_389646 ; 
   reg __389646_389646;
   reg _389647_389647 ; 
   reg __389647_389647;
   reg _389648_389648 ; 
   reg __389648_389648;
   reg _389649_389649 ; 
   reg __389649_389649;
   reg _389650_389650 ; 
   reg __389650_389650;
   reg _389651_389651 ; 
   reg __389651_389651;
   reg _389652_389652 ; 
   reg __389652_389652;
   reg _389653_389653 ; 
   reg __389653_389653;
   reg _389654_389654 ; 
   reg __389654_389654;
   reg _389655_389655 ; 
   reg __389655_389655;
   reg _389656_389656 ; 
   reg __389656_389656;
   reg _389657_389657 ; 
   reg __389657_389657;
   reg _389658_389658 ; 
   reg __389658_389658;
   reg _389659_389659 ; 
   reg __389659_389659;
   reg _389660_389660 ; 
   reg __389660_389660;
   reg _389661_389661 ; 
   reg __389661_389661;
   reg _389662_389662 ; 
   reg __389662_389662;
   reg _389663_389663 ; 
   reg __389663_389663;
   reg _389664_389664 ; 
   reg __389664_389664;
   reg _389665_389665 ; 
   reg __389665_389665;
   reg _389666_389666 ; 
   reg __389666_389666;
   reg _389667_389667 ; 
   reg __389667_389667;
   reg _389668_389668 ; 
   reg __389668_389668;
   reg _389669_389669 ; 
   reg __389669_389669;
   reg _389670_389670 ; 
   reg __389670_389670;
   reg _389671_389671 ; 
   reg __389671_389671;
   reg _389672_389672 ; 
   reg __389672_389672;
   reg _389673_389673 ; 
   reg __389673_389673;
   reg _389674_389674 ; 
   reg __389674_389674;
   reg _389675_389675 ; 
   reg __389675_389675;
   reg _389676_389676 ; 
   reg __389676_389676;
   reg _389677_389677 ; 
   reg __389677_389677;
   reg _389678_389678 ; 
   reg __389678_389678;
   reg _389679_389679 ; 
   reg __389679_389679;
   reg _389680_389680 ; 
   reg __389680_389680;
   reg _389681_389681 ; 
   reg __389681_389681;
   reg _389682_389682 ; 
   reg __389682_389682;
   reg _389683_389683 ; 
   reg __389683_389683;
   reg _389684_389684 ; 
   reg __389684_389684;
   reg _389685_389685 ; 
   reg __389685_389685;
   reg _389686_389686 ; 
   reg __389686_389686;
   reg _389687_389687 ; 
   reg __389687_389687;
   reg _389688_389688 ; 
   reg __389688_389688;
   reg _389689_389689 ; 
   reg __389689_389689;
   reg _389690_389690 ; 
   reg __389690_389690;
   reg _389691_389691 ; 
   reg __389691_389691;
   reg _389692_389692 ; 
   reg __389692_389692;
   reg _389693_389693 ; 
   reg __389693_389693;
   reg _389694_389694 ; 
   reg __389694_389694;
   reg _389695_389695 ; 
   reg __389695_389695;
   reg _389696_389696 ; 
   reg __389696_389696;
   reg _389697_389697 ; 
   reg __389697_389697;
   reg _389698_389698 ; 
   reg __389698_389698;
   reg _389699_389699 ; 
   reg __389699_389699;
   reg _389700_389700 ; 
   reg __389700_389700;
   reg _389701_389701 ; 
   reg __389701_389701;
   reg _389702_389702 ; 
   reg __389702_389702;
   reg _389703_389703 ; 
   reg __389703_389703;
   reg _389704_389704 ; 
   reg __389704_389704;
   reg _389705_389705 ; 
   reg __389705_389705;
   reg _389706_389706 ; 
   reg __389706_389706;
   reg _389707_389707 ; 
   reg __389707_389707;
   reg _389708_389708 ; 
   reg __389708_389708;
   reg _389709_389709 ; 
   reg __389709_389709;
   reg _389710_389710 ; 
   reg __389710_389710;
   reg _389711_389711 ; 
   reg __389711_389711;
   reg _389712_389712 ; 
   reg __389712_389712;
   reg _389713_389713 ; 
   reg __389713_389713;
   reg _389714_389714 ; 
   reg __389714_389714;
   reg _389715_389715 ; 
   reg __389715_389715;
   reg _389716_389716 ; 
   reg __389716_389716;
   reg _389717_389717 ; 
   reg __389717_389717;
   reg _389718_389718 ; 
   reg __389718_389718;
   reg _389719_389719 ; 
   reg __389719_389719;
   reg _389720_389720 ; 
   reg __389720_389720;
   reg _389721_389721 ; 
   reg __389721_389721;
   reg _389722_389722 ; 
   reg __389722_389722;
   reg _389723_389723 ; 
   reg __389723_389723;
   reg _389724_389724 ; 
   reg __389724_389724;
   reg _389725_389725 ; 
   reg __389725_389725;
   reg _389726_389726 ; 
   reg __389726_389726;
   reg _389727_389727 ; 
   reg __389727_389727;
   reg _389728_389728 ; 
   reg __389728_389728;
   reg _389729_389729 ; 
   reg __389729_389729;
   reg _389730_389730 ; 
   reg __389730_389730;
   reg _389731_389731 ; 
   reg __389731_389731;
   reg _389732_389732 ; 
   reg __389732_389732;
   reg _389733_389733 ; 
   reg __389733_389733;
   reg _389734_389734 ; 
   reg __389734_389734;
   reg _389735_389735 ; 
   reg __389735_389735;
   reg _389736_389736 ; 
   reg __389736_389736;
   reg _389737_389737 ; 
   reg __389737_389737;
   reg _389738_389738 ; 
   reg __389738_389738;
   reg _389739_389739 ; 
   reg __389739_389739;
   reg _389740_389740 ; 
   reg __389740_389740;
   reg _389741_389741 ; 
   reg __389741_389741;
   reg _389742_389742 ; 
   reg __389742_389742;
   reg _389743_389743 ; 
   reg __389743_389743;
   reg _389744_389744 ; 
   reg __389744_389744;
   reg _389745_389745 ; 
   reg __389745_389745;
   reg _389746_389746 ; 
   reg __389746_389746;
   reg _389747_389747 ; 
   reg __389747_389747;
   reg _389748_389748 ; 
   reg __389748_389748;
   reg _389749_389749 ; 
   reg __389749_389749;
   reg _389750_389750 ; 
   reg __389750_389750;
   reg _389751_389751 ; 
   reg __389751_389751;
   reg _389752_389752 ; 
   reg __389752_389752;
   reg _389753_389753 ; 
   reg __389753_389753;
   reg _389754_389754 ; 
   reg __389754_389754;
   reg _389755_389755 ; 
   reg __389755_389755;
   reg _389756_389756 ; 
   reg __389756_389756;
   reg _389757_389757 ; 
   reg __389757_389757;
   reg _389758_389758 ; 
   reg __389758_389758;
   reg _389759_389759 ; 
   reg __389759_389759;
   reg _389760_389760 ; 
   reg __389760_389760;
   reg _389761_389761 ; 
   reg __389761_389761;
   reg _389762_389762 ; 
   reg __389762_389762;
   reg _389763_389763 ; 
   reg __389763_389763;
   reg _389764_389764 ; 
   reg __389764_389764;
   reg _389765_389765 ; 
   reg __389765_389765;
   reg _389766_389766 ; 
   reg __389766_389766;
   reg _389767_389767 ; 
   reg __389767_389767;
   reg _389768_389768 ; 
   reg __389768_389768;
   reg _389769_389769 ; 
   reg __389769_389769;
   reg _389770_389770 ; 
   reg __389770_389770;
   reg _389771_389771 ; 
   reg __389771_389771;
   reg _389772_389772 ; 
   reg __389772_389772;
   reg _389773_389773 ; 
   reg __389773_389773;
   reg _389774_389774 ; 
   reg __389774_389774;
   reg _389775_389775 ; 
   reg __389775_389775;
   reg _389776_389776 ; 
   reg __389776_389776;
   reg _389777_389777 ; 
   reg __389777_389777;
   reg _389778_389778 ; 
   reg __389778_389778;
   reg _389779_389779 ; 
   reg __389779_389779;
   reg _389780_389780 ; 
   reg __389780_389780;
   reg _389781_389781 ; 
   reg __389781_389781;
   reg _389782_389782 ; 
   reg __389782_389782;
   reg _389783_389783 ; 
   reg __389783_389783;
   reg _389784_389784 ; 
   reg __389784_389784;
   reg _389785_389785 ; 
   reg __389785_389785;
   reg _389786_389786 ; 
   reg __389786_389786;
   reg _389787_389787 ; 
   reg __389787_389787;
   reg _389788_389788 ; 
   reg __389788_389788;
   reg _389789_389789 ; 
   reg __389789_389789;
   reg _389790_389790 ; 
   reg __389790_389790;
   reg _389791_389791 ; 
   reg __389791_389791;
   reg _389792_389792 ; 
   reg __389792_389792;
   reg _389793_389793 ; 
   reg __389793_389793;
   reg _389794_389794 ; 
   reg __389794_389794;
   reg _389795_389795 ; 
   reg __389795_389795;
   reg _389796_389796 ; 
   reg __389796_389796;
   reg _389797_389797 ; 
   reg __389797_389797;
   reg _389798_389798 ; 
   reg __389798_389798;
   reg _389799_389799 ; 
   reg __389799_389799;
   reg _389800_389800 ; 
   reg __389800_389800;
   reg _389801_389801 ; 
   reg __389801_389801;
   reg _389802_389802 ; 
   reg __389802_389802;
   reg _389803_389803 ; 
   reg __389803_389803;
   reg _389804_389804 ; 
   reg __389804_389804;
   reg _389805_389805 ; 
   reg __389805_389805;
   reg _389806_389806 ; 
   reg __389806_389806;
   reg _389807_389807 ; 
   reg __389807_389807;
   reg _389808_389808 ; 
   reg __389808_389808;
   reg _389809_389809 ; 
   reg __389809_389809;
   reg _389810_389810 ; 
   reg __389810_389810;
   reg _389811_389811 ; 
   reg __389811_389811;
   reg _389812_389812 ; 
   reg __389812_389812;
   reg _389813_389813 ; 
   reg __389813_389813;
   reg _389814_389814 ; 
   reg __389814_389814;
   reg _389815_389815 ; 
   reg __389815_389815;
   reg _389816_389816 ; 
   reg __389816_389816;
   reg _389817_389817 ; 
   reg __389817_389817;
   reg _389818_389818 ; 
   reg __389818_389818;
   reg _389819_389819 ; 
   reg __389819_389819;
   reg _389820_389820 ; 
   reg __389820_389820;
   reg _389821_389821 ; 
   reg __389821_389821;
   reg _389822_389822 ; 
   reg __389822_389822;
   reg _389823_389823 ; 
   reg __389823_389823;
   reg _389824_389824 ; 
   reg __389824_389824;
   reg _389825_389825 ; 
   reg __389825_389825;
   reg _389826_389826 ; 
   reg __389826_389826;
   reg _389827_389827 ; 
   reg __389827_389827;
   reg _389828_389828 ; 
   reg __389828_389828;
   reg _389829_389829 ; 
   reg __389829_389829;
   reg _389830_389830 ; 
   reg __389830_389830;
   reg _389831_389831 ; 
   reg __389831_389831;
   reg _389832_389832 ; 
   reg __389832_389832;
   reg _389833_389833 ; 
   reg __389833_389833;
   reg _389834_389834 ; 
   reg __389834_389834;
   reg _389835_389835 ; 
   reg __389835_389835;
   reg _389836_389836 ; 
   reg __389836_389836;
   reg _389837_389837 ; 
   reg __389837_389837;
   reg _389838_389838 ; 
   reg __389838_389838;
   reg _389839_389839 ; 
   reg __389839_389839;
   reg _389840_389840 ; 
   reg __389840_389840;
   reg _389841_389841 ; 
   reg __389841_389841;
   reg _389842_389842 ; 
   reg __389842_389842;
   reg _389843_389843 ; 
   reg __389843_389843;
   reg _389844_389844 ; 
   reg __389844_389844;
   reg _389845_389845 ; 
   reg __389845_389845;
   reg _389846_389846 ; 
   reg __389846_389846;
   reg _389847_389847 ; 
   reg __389847_389847;
   reg _389848_389848 ; 
   reg __389848_389848;
   reg _389849_389849 ; 
   reg __389849_389849;
   reg _389850_389850 ; 
   reg __389850_389850;
   reg _389851_389851 ; 
   reg __389851_389851;
   reg _389852_389852 ; 
   reg __389852_389852;
   reg _389853_389853 ; 
   reg __389853_389853;
   reg _389854_389854 ; 
   reg __389854_389854;
   reg _389855_389855 ; 
   reg __389855_389855;
   reg _389856_389856 ; 
   reg __389856_389856;
   reg _389857_389857 ; 
   reg __389857_389857;
   reg _389858_389858 ; 
   reg __389858_389858;
   reg _389859_389859 ; 
   reg __389859_389859;
   reg _389860_389860 ; 
   reg __389860_389860;
   reg _389861_389861 ; 
   reg __389861_389861;
   reg _389862_389862 ; 
   reg __389862_389862;
   reg _389863_389863 ; 
   reg __389863_389863;
   reg _389864_389864 ; 
   reg __389864_389864;
   reg _389865_389865 ; 
   reg __389865_389865;
   reg _389866_389866 ; 
   reg __389866_389866;
   reg _389867_389867 ; 
   reg __389867_389867;
   reg _389868_389868 ; 
   reg __389868_389868;
   reg _389869_389869 ; 
   reg __389869_389869;
   reg _389870_389870 ; 
   reg __389870_389870;
   reg _389871_389871 ; 
   reg __389871_389871;
   reg _389872_389872 ; 
   reg __389872_389872;
   reg _389873_389873 ; 
   reg __389873_389873;
   reg _389874_389874 ; 
   reg __389874_389874;
   reg _389875_389875 ; 
   reg __389875_389875;
   reg _389876_389876 ; 
   reg __389876_389876;
   reg _389877_389877 ; 
   reg __389877_389877;
   reg _389878_389878 ; 
   reg __389878_389878;
   reg _389879_389879 ; 
   reg __389879_389879;
   reg _389880_389880 ; 
   reg __389880_389880;
   reg _389881_389881 ; 
   reg __389881_389881;
   reg _389882_389882 ; 
   reg __389882_389882;
   reg _389883_389883 ; 
   reg __389883_389883;
   reg _389884_389884 ; 
   reg __389884_389884;
   reg _389885_389885 ; 
   reg __389885_389885;
   reg _389886_389886 ; 
   reg __389886_389886;
   reg _389887_389887 ; 
   reg __389887_389887;
   reg _389888_389888 ; 
   reg __389888_389888;
   reg _389889_389889 ; 
   reg __389889_389889;
   reg _389890_389890 ; 
   reg __389890_389890;
   reg _389891_389891 ; 
   reg __389891_389891;
   reg _389892_389892 ; 
   reg __389892_389892;
   reg _389893_389893 ; 
   reg __389893_389893;
   reg _389894_389894 ; 
   reg __389894_389894;
   reg _389895_389895 ; 
   reg __389895_389895;
   reg _389896_389896 ; 
   reg __389896_389896;
   reg _389897_389897 ; 
   reg __389897_389897;
   reg _389898_389898 ; 
   reg __389898_389898;
   reg _389899_389899 ; 
   reg __389899_389899;
   reg _389900_389900 ; 
   reg __389900_389900;
   reg _389901_389901 ; 
   reg __389901_389901;
   reg _389902_389902 ; 
   reg __389902_389902;
   reg _389903_389903 ; 
   reg __389903_389903;
   reg _389904_389904 ; 
   reg __389904_389904;
   reg _389905_389905 ; 
   reg __389905_389905;
   reg _389906_389906 ; 
   reg __389906_389906;
   reg _389907_389907 ; 
   reg __389907_389907;
   reg _389908_389908 ; 
   reg __389908_389908;
   reg _389909_389909 ; 
   reg __389909_389909;
   reg _389910_389910 ; 
   reg __389910_389910;
   reg _389911_389911 ; 
   reg __389911_389911;
   reg _389912_389912 ; 
   reg __389912_389912;
   reg _389913_389913 ; 
   reg __389913_389913;
   reg _389914_389914 ; 
   reg __389914_389914;
   reg _389915_389915 ; 
   reg __389915_389915;
   reg _389916_389916 ; 
   reg __389916_389916;
   reg _389917_389917 ; 
   reg __389917_389917;
   reg _389918_389918 ; 
   reg __389918_389918;
   reg _389919_389919 ; 
   reg __389919_389919;
   reg _389920_389920 ; 
   reg __389920_389920;
   reg _389921_389921 ; 
   reg __389921_389921;
   reg _389922_389922 ; 
   reg __389922_389922;
   reg _389923_389923 ; 
   reg __389923_389923;
   reg _389924_389924 ; 
   reg __389924_389924;
   reg _389925_389925 ; 
   reg __389925_389925;
   reg _389926_389926 ; 
   reg __389926_389926;
   reg _389927_389927 ; 
   reg __389927_389927;
   reg _389928_389928 ; 
   reg __389928_389928;
   reg _389929_389929 ; 
   reg __389929_389929;
   reg _389930_389930 ; 
   reg __389930_389930;
   reg _389931_389931 ; 
   reg __389931_389931;
   reg _389932_389932 ; 
   reg __389932_389932;
   reg _389933_389933 ; 
   reg __389933_389933;
   reg _389934_389934 ; 
   reg __389934_389934;
   reg _389935_389935 ; 
   reg __389935_389935;
   reg _389936_389936 ; 
   reg __389936_389936;
   reg _389937_389937 ; 
   reg __389937_389937;
   reg _389938_389938 ; 
   reg __389938_389938;
   reg _389939_389939 ; 
   reg __389939_389939;
   reg _389940_389940 ; 
   reg __389940_389940;
   reg _389941_389941 ; 
   reg __389941_389941;
   reg _389942_389942 ; 
   reg __389942_389942;
   reg _389943_389943 ; 
   reg __389943_389943;
   reg _389944_389944 ; 
   reg __389944_389944;
   reg _389945_389945 ; 
   reg __389945_389945;
   reg _389946_389946 ; 
   reg __389946_389946;
   reg _389947_389947 ; 
   reg __389947_389947;
   reg _389948_389948 ; 
   reg __389948_389948;
   reg _389949_389949 ; 
   reg __389949_389949;
   reg _389950_389950 ; 
   reg __389950_389950;
   reg _389951_389951 ; 
   reg __389951_389951;
   reg _389952_389952 ; 
   reg __389952_389952;
   reg _389953_389953 ; 
   reg __389953_389953;
   reg _389954_389954 ; 
   reg __389954_389954;
   reg _389955_389955 ; 
   reg __389955_389955;
   reg _389956_389956 ; 
   reg __389956_389956;
   reg _389957_389957 ; 
   reg __389957_389957;
   reg _389958_389958 ; 
   reg __389958_389958;
   reg _389959_389959 ; 
   reg __389959_389959;
   reg _389960_389960 ; 
   reg __389960_389960;
   reg _389961_389961 ; 
   reg __389961_389961;
   reg _389962_389962 ; 
   reg __389962_389962;
   reg _389963_389963 ; 
   reg __389963_389963;
   reg _389964_389964 ; 
   reg __389964_389964;
   reg _389965_389965 ; 
   reg __389965_389965;
   reg _389966_389966 ; 
   reg __389966_389966;
   reg _389967_389967 ; 
   reg __389967_389967;
   reg _389968_389968 ; 
   reg __389968_389968;
   reg _389969_389969 ; 
   reg __389969_389969;
   reg _389970_389970 ; 
   reg __389970_389970;
   reg _389971_389971 ; 
   reg __389971_389971;
   reg _389972_389972 ; 
   reg __389972_389972;
   reg _389973_389973 ; 
   reg __389973_389973;
   reg _389974_389974 ; 
   reg __389974_389974;
   reg _389975_389975 ; 
   reg __389975_389975;
   reg _389976_389976 ; 
   reg __389976_389976;
   reg _389977_389977 ; 
   reg __389977_389977;
   reg _389978_389978 ; 
   reg __389978_389978;
   reg _389979_389979 ; 
   reg __389979_389979;
   reg _389980_389980 ; 
   reg __389980_389980;
   reg _389981_389981 ; 
   reg __389981_389981;
   reg _389982_389982 ; 
   reg __389982_389982;
   reg _389983_389983 ; 
   reg __389983_389983;
   reg _389984_389984 ; 
   reg __389984_389984;
   reg _389985_389985 ; 
   reg __389985_389985;
   reg _389986_389986 ; 
   reg __389986_389986;
   reg _389987_389987 ; 
   reg __389987_389987;
   reg _389988_389988 ; 
   reg __389988_389988;
   reg _389989_389989 ; 
   reg __389989_389989;
   reg _389990_389990 ; 
   reg __389990_389990;
   reg _389991_389991 ; 
   reg __389991_389991;
   reg _389992_389992 ; 
   reg __389992_389992;
   reg _389993_389993 ; 
   reg __389993_389993;
   reg _389994_389994 ; 
   reg __389994_389994;
   reg _389995_389995 ; 
   reg __389995_389995;
   reg _389996_389996 ; 
   reg __389996_389996;
   reg _389997_389997 ; 
   reg __389997_389997;
   reg _389998_389998 ; 
   reg __389998_389998;
   reg _389999_389999 ; 
   reg __389999_389999;
   reg _390000_390000 ; 
   reg __390000_390000;
   reg _390001_390001 ; 
   reg __390001_390001;
   reg _390002_390002 ; 
   reg __390002_390002;
   reg _390003_390003 ; 
   reg __390003_390003;
   reg _390004_390004 ; 
   reg __390004_390004;
   reg _390005_390005 ; 
   reg __390005_390005;
   reg _390006_390006 ; 
   reg __390006_390006;
   reg _390007_390007 ; 
   reg __390007_390007;
   reg _390008_390008 ; 
   reg __390008_390008;
   reg _390009_390009 ; 
   reg __390009_390009;
   reg _390010_390010 ; 
   reg __390010_390010;
   reg _390011_390011 ; 
   reg __390011_390011;
   reg _390012_390012 ; 
   reg __390012_390012;
   reg _390013_390013 ; 
   reg __390013_390013;
   reg _390014_390014 ; 
   reg __390014_390014;
   reg _390015_390015 ; 
   reg __390015_390015;
   reg _390016_390016 ; 
   reg __390016_390016;
   reg _390017_390017 ; 
   reg __390017_390017;
   reg _390018_390018 ; 
   reg __390018_390018;
   reg _390019_390019 ; 
   reg __390019_390019;
   reg _390020_390020 ; 
   reg __390020_390020;
   reg _390021_390021 ; 
   reg __390021_390021;
   reg _390022_390022 ; 
   reg __390022_390022;
   reg _390023_390023 ; 
   reg __390023_390023;
   reg _390024_390024 ; 
   reg __390024_390024;
   reg _390025_390025 ; 
   reg __390025_390025;
   reg _390026_390026 ; 
   reg __390026_390026;
   reg _390027_390027 ; 
   reg __390027_390027;
   reg _390028_390028 ; 
   reg __390028_390028;
   reg _390029_390029 ; 
   reg __390029_390029;
   reg _390030_390030 ; 
   reg __390030_390030;
   reg _390031_390031 ; 
   reg __390031_390031;
   reg _390032_390032 ; 
   reg __390032_390032;
   reg _390033_390033 ; 
   reg __390033_390033;
   reg _390034_390034 ; 
   reg __390034_390034;
   reg _390035_390035 ; 
   reg __390035_390035;
   reg _390036_390036 ; 
   reg __390036_390036;
   reg _390037_390037 ; 
   reg __390037_390037;
   reg _390038_390038 ; 
   reg __390038_390038;
   reg _390039_390039 ; 
   reg __390039_390039;
   reg _390040_390040 ; 
   reg __390040_390040;
   reg _390041_390041 ; 
   reg __390041_390041;
   reg _390042_390042 ; 
   reg __390042_390042;
   reg _390043_390043 ; 
   reg __390043_390043;
   reg _390044_390044 ; 
   reg __390044_390044;
   reg _390045_390045 ; 
   reg __390045_390045;
   reg _390046_390046 ; 
   reg __390046_390046;
   reg _390047_390047 ; 
   reg __390047_390047;
   reg _390048_390048 ; 
   reg __390048_390048;
   reg _390049_390049 ; 
   reg __390049_390049;
   reg _390050_390050 ; 
   reg __390050_390050;
   reg _390051_390051 ; 
   reg __390051_390051;
   reg _390052_390052 ; 
   reg __390052_390052;
   reg _390053_390053 ; 
   reg __390053_390053;
   reg _390054_390054 ; 
   reg __390054_390054;
   reg _390055_390055 ; 
   reg __390055_390055;
   reg _390056_390056 ; 
   reg __390056_390056;
   reg _390057_390057 ; 
   reg __390057_390057;
   reg _390058_390058 ; 
   reg __390058_390058;
   reg _390059_390059 ; 
   reg __390059_390059;
   reg _390060_390060 ; 
   reg __390060_390060;
   reg _390061_390061 ; 
   reg __390061_390061;
   reg _390062_390062 ; 
   reg __390062_390062;
   reg _390063_390063 ; 
   reg __390063_390063;
   reg _390064_390064 ; 
   reg __390064_390064;
   reg _390065_390065 ; 
   reg __390065_390065;
   reg _390066_390066 ; 
   reg __390066_390066;
   reg _390067_390067 ; 
   reg __390067_390067;
   reg _390068_390068 ; 
   reg __390068_390068;
   reg _390069_390069 ; 
   reg __390069_390069;
   reg _390070_390070 ; 
   reg __390070_390070;
   reg _390071_390071 ; 
   reg __390071_390071;
   reg _390072_390072 ; 
   reg __390072_390072;
   reg _390073_390073 ; 
   reg __390073_390073;
   reg _390074_390074 ; 
   reg __390074_390074;
   reg _390075_390075 ; 
   reg __390075_390075;
   reg _390076_390076 ; 
   reg __390076_390076;
   reg _390077_390077 ; 
   reg __390077_390077;
   reg _390078_390078 ; 
   reg __390078_390078;
   reg _390079_390079 ; 
   reg __390079_390079;
   reg _390080_390080 ; 
   reg __390080_390080;
   reg _390081_390081 ; 
   reg __390081_390081;
   reg _390082_390082 ; 
   reg __390082_390082;
   reg _390083_390083 ; 
   reg __390083_390083;
   reg _390084_390084 ; 
   reg __390084_390084;
   reg _390085_390085 ; 
   reg __390085_390085;
   reg _390086_390086 ; 
   reg __390086_390086;
   reg _390087_390087 ; 
   reg __390087_390087;
   reg _390088_390088 ; 
   reg __390088_390088;
   reg _390089_390089 ; 
   reg __390089_390089;
   reg _390090_390090 ; 
   reg __390090_390090;
   reg _390091_390091 ; 
   reg __390091_390091;
   reg _390092_390092 ; 
   reg __390092_390092;
   reg _390093_390093 ; 
   reg __390093_390093;
   reg _390094_390094 ; 
   reg __390094_390094;
   reg _390095_390095 ; 
   reg __390095_390095;
   reg _390096_390096 ; 
   reg __390096_390096;
   reg _390097_390097 ; 
   reg __390097_390097;
   reg _390098_390098 ; 
   reg __390098_390098;
   reg _390099_390099 ; 
   reg __390099_390099;
   reg _390100_390100 ; 
   reg __390100_390100;
   reg _390101_390101 ; 
   reg __390101_390101;
   reg _390102_390102 ; 
   reg __390102_390102;
   reg _390103_390103 ; 
   reg __390103_390103;
   reg _390104_390104 ; 
   reg __390104_390104;
   reg _390105_390105 ; 
   reg __390105_390105;
   reg _390106_390106 ; 
   reg __390106_390106;
   reg _390107_390107 ; 
   reg __390107_390107;
   reg _390108_390108 ; 
   reg __390108_390108;
   reg _390109_390109 ; 
   reg __390109_390109;
   reg _390110_390110 ; 
   reg __390110_390110;
   reg _390111_390111 ; 
   reg __390111_390111;
   reg _390112_390112 ; 
   reg __390112_390112;
   reg _390113_390113 ; 
   reg __390113_390113;
   reg _390114_390114 ; 
   reg __390114_390114;
   reg _390115_390115 ; 
   reg __390115_390115;
   reg _390116_390116 ; 
   reg __390116_390116;
   reg _390117_390117 ; 
   reg __390117_390117;
   reg _390118_390118 ; 
   reg __390118_390118;
   reg _390119_390119 ; 
   reg __390119_390119;
   reg _390120_390120 ; 
   reg __390120_390120;
   reg _390121_390121 ; 
   reg __390121_390121;
   reg _390122_390122 ; 
   reg __390122_390122;
   reg _390123_390123 ; 
   reg __390123_390123;
   reg _390124_390124 ; 
   reg __390124_390124;
   reg _390125_390125 ; 
   reg __390125_390125;
   reg _390126_390126 ; 
   reg __390126_390126;
   reg _390127_390127 ; 
   reg __390127_390127;
   reg _390128_390128 ; 
   reg __390128_390128;
   reg _390129_390129 ; 
   reg __390129_390129;
   reg _390130_390130 ; 
   reg __390130_390130;
   reg _390131_390131 ; 
   reg __390131_390131;
   reg _390132_390132 ; 
   reg __390132_390132;
   reg _390133_390133 ; 
   reg __390133_390133;
   reg _390134_390134 ; 
   reg __390134_390134;
   reg _390135_390135 ; 
   reg __390135_390135;
   reg _390136_390136 ; 
   reg __390136_390136;
   reg _390137_390137 ; 
   reg __390137_390137;
   reg _390138_390138 ; 
   reg __390138_390138;
   reg _390139_390139 ; 
   reg __390139_390139;
   reg _390140_390140 ; 
   reg __390140_390140;
   reg _390141_390141 ; 
   reg __390141_390141;
   reg _390142_390142 ; 
   reg __390142_390142;
   reg _390143_390143 ; 
   reg __390143_390143;
   reg _390144_390144 ; 
   reg __390144_390144;
   reg _390145_390145 ; 
   reg __390145_390145;
   reg _390146_390146 ; 
   reg __390146_390146;
   reg _390147_390147 ; 
   reg __390147_390147;
   reg _390148_390148 ; 
   reg __390148_390148;
   reg _390149_390149 ; 
   reg __390149_390149;
   reg _390150_390150 ; 
   reg __390150_390150;
   reg _390151_390151 ; 
   reg __390151_390151;
   reg _390152_390152 ; 
   reg __390152_390152;
   reg _390153_390153 ; 
   reg __390153_390153;
   reg _390154_390154 ; 
   reg __390154_390154;
   reg _390155_390155 ; 
   reg __390155_390155;
   reg _390156_390156 ; 
   reg __390156_390156;
   reg _390157_390157 ; 
   reg __390157_390157;
   reg _390158_390158 ; 
   reg __390158_390158;
   reg _390159_390159 ; 
   reg __390159_390159;
   reg _390160_390160 ; 
   reg __390160_390160;
   reg _390161_390161 ; 
   reg __390161_390161;
   reg _390162_390162 ; 
   reg __390162_390162;
   reg _390163_390163 ; 
   reg __390163_390163;
   reg _390164_390164 ; 
   reg __390164_390164;
   reg _390165_390165 ; 
   reg __390165_390165;
   reg _390166_390166 ; 
   reg __390166_390166;
   reg _390167_390167 ; 
   reg __390167_390167;
   reg _390168_390168 ; 
   reg __390168_390168;
   reg _390169_390169 ; 
   reg __390169_390169;
   reg _390170_390170 ; 
   reg __390170_390170;
   reg _390171_390171 ; 
   reg __390171_390171;
   reg _390172_390172 ; 
   reg __390172_390172;
   reg _390173_390173 ; 
   reg __390173_390173;
   reg _390174_390174 ; 
   reg __390174_390174;
   reg _390175_390175 ; 
   reg __390175_390175;
   reg _390176_390176 ; 
   reg __390176_390176;
   reg _390177_390177 ; 
   reg __390177_390177;
   reg _390178_390178 ; 
   reg __390178_390178;
   reg _390179_390179 ; 
   reg __390179_390179;
   reg _390180_390180 ; 
   reg __390180_390180;
   reg _390181_390181 ; 
   reg __390181_390181;
   reg _390182_390182 ; 
   reg __390182_390182;
   reg _390183_390183 ; 
   reg __390183_390183;
   reg _390184_390184 ; 
   reg __390184_390184;
   reg _390185_390185 ; 
   reg __390185_390185;
   reg _390186_390186 ; 
   reg __390186_390186;
   reg _390187_390187 ; 
   reg __390187_390187;
   reg _390188_390188 ; 
   reg __390188_390188;
   reg _390189_390189 ; 
   reg __390189_390189;
   reg _390190_390190 ; 
   reg __390190_390190;
   reg _390191_390191 ; 
   reg __390191_390191;
   reg _390192_390192 ; 
   reg __390192_390192;
   reg _390193_390193 ; 
   reg __390193_390193;
   reg _390194_390194 ; 
   reg __390194_390194;
   reg _390195_390195 ; 
   reg __390195_390195;
   reg _390196_390196 ; 
   reg __390196_390196;
   reg _390197_390197 ; 
   reg __390197_390197;
   reg _390198_390198 ; 
   reg __390198_390198;
   reg _390199_390199 ; 
   reg __390199_390199;
   reg _390200_390200 ; 
   reg __390200_390200;
   reg _390201_390201 ; 
   reg __390201_390201;
   reg _390202_390202 ; 
   reg __390202_390202;
   reg _390203_390203 ; 
   reg __390203_390203;
   reg _390204_390204 ; 
   reg __390204_390204;
   reg _390205_390205 ; 
   reg __390205_390205;
   reg _390206_390206 ; 
   reg __390206_390206;
   reg _390207_390207 ; 
   reg __390207_390207;
   reg _390208_390208 ; 
   reg __390208_390208;
   reg _390209_390209 ; 
   reg __390209_390209;
   reg _390210_390210 ; 
   reg __390210_390210;
   reg _390211_390211 ; 
   reg __390211_390211;
   reg _390212_390212 ; 
   reg __390212_390212;
   reg _390213_390213 ; 
   reg __390213_390213;
   reg _390214_390214 ; 
   reg __390214_390214;
   reg _390215_390215 ; 
   reg __390215_390215;
   reg _390216_390216 ; 
   reg __390216_390216;
   reg _390217_390217 ; 
   reg __390217_390217;
   reg _390218_390218 ; 
   reg __390218_390218;
   reg _390219_390219 ; 
   reg __390219_390219;
   reg _390220_390220 ; 
   reg __390220_390220;
   reg _390221_390221 ; 
   reg __390221_390221;
   reg _390222_390222 ; 
   reg __390222_390222;
   reg _390223_390223 ; 
   reg __390223_390223;
   reg _390224_390224 ; 
   reg __390224_390224;
   reg _390225_390225 ; 
   reg __390225_390225;
   reg _390226_390226 ; 
   reg __390226_390226;
   reg _390227_390227 ; 
   reg __390227_390227;
   reg _390228_390228 ; 
   reg __390228_390228;
   reg _390229_390229 ; 
   reg __390229_390229;
   reg _390230_390230 ; 
   reg __390230_390230;
   reg _390231_390231 ; 
   reg __390231_390231;
   reg _390232_390232 ; 
   reg __390232_390232;
   reg _390233_390233 ; 
   reg __390233_390233;
   reg _390234_390234 ; 
   reg __390234_390234;
   reg _390235_390235 ; 
   reg __390235_390235;
   reg _390236_390236 ; 
   reg __390236_390236;
   reg _390237_390237 ; 
   reg __390237_390237;
   reg _390238_390238 ; 
   reg __390238_390238;
   reg _390239_390239 ; 
   reg __390239_390239;
   reg _390240_390240 ; 
   reg __390240_390240;
   reg _390241_390241 ; 
   reg __390241_390241;
   reg _390242_390242 ; 
   reg __390242_390242;
   reg _390243_390243 ; 
   reg __390243_390243;
   reg _390244_390244 ; 
   reg __390244_390244;
   reg _390245_390245 ; 
   reg __390245_390245;
   reg _390246_390246 ; 
   reg __390246_390246;
   reg _390247_390247 ; 
   reg __390247_390247;
   reg _390248_390248 ; 
   reg __390248_390248;
   reg _390249_390249 ; 
   reg __390249_390249;
   reg _390250_390250 ; 
   reg __390250_390250;
   reg _390251_390251 ; 
   reg __390251_390251;
   reg _390252_390252 ; 
   reg __390252_390252;
   reg _390253_390253 ; 
   reg __390253_390253;
   reg _390254_390254 ; 
   reg __390254_390254;
   reg _390255_390255 ; 
   reg __390255_390255;
   reg _390256_390256 ; 
   reg __390256_390256;
   reg _390257_390257 ; 
   reg __390257_390257;
   reg _390258_390258 ; 
   reg __390258_390258;
   reg _390259_390259 ; 
   reg __390259_390259;
   reg _390260_390260 ; 
   reg __390260_390260;
   reg _390261_390261 ; 
   reg __390261_390261;
   reg _390262_390262 ; 
   reg __390262_390262;
   reg _390263_390263 ; 
   reg __390263_390263;
   reg _390264_390264 ; 
   reg __390264_390264;
   reg _390265_390265 ; 
   reg __390265_390265;
   reg _390266_390266 ; 
   reg __390266_390266;
   reg _390267_390267 ; 
   reg __390267_390267;
   reg _390268_390268 ; 
   reg __390268_390268;
   reg _390269_390269 ; 
   reg __390269_390269;
   reg _390270_390270 ; 
   reg __390270_390270;
   reg _390271_390271 ; 
   reg __390271_390271;
   reg _390272_390272 ; 
   reg __390272_390272;
   reg _390273_390273 ; 
   reg __390273_390273;
   reg _390274_390274 ; 
   reg __390274_390274;
   reg _390275_390275 ; 
   reg __390275_390275;
   reg _390276_390276 ; 
   reg __390276_390276;
   reg _390277_390277 ; 
   reg __390277_390277;
   reg _390278_390278 ; 
   reg __390278_390278;
   reg _390279_390279 ; 
   reg __390279_390279;
   reg _390280_390280 ; 
   reg __390280_390280;
   reg _390281_390281 ; 
   reg __390281_390281;
   reg _390282_390282 ; 
   reg __390282_390282;
   reg _390283_390283 ; 
   reg __390283_390283;
   reg _390284_390284 ; 
   reg __390284_390284;
   reg _390285_390285 ; 
   reg __390285_390285;
   reg _390286_390286 ; 
   reg __390286_390286;
   reg _390287_390287 ; 
   reg __390287_390287;
   reg _390288_390288 ; 
   reg __390288_390288;
   reg _390289_390289 ; 
   reg __390289_390289;
   reg _390290_390290 ; 
   reg __390290_390290;
   reg _390291_390291 ; 
   reg __390291_390291;
   reg _390292_390292 ; 
   reg __390292_390292;
   reg _390293_390293 ; 
   reg __390293_390293;
   reg _390294_390294 ; 
   reg __390294_390294;
   reg _390295_390295 ; 
   reg __390295_390295;
   reg _390296_390296 ; 
   reg __390296_390296;
   reg _390297_390297 ; 
   reg __390297_390297;
   reg _390298_390298 ; 
   reg __390298_390298;
   reg _390299_390299 ; 
   reg __390299_390299;
   reg _390300_390300 ; 
   reg __390300_390300;
   reg _390301_390301 ; 
   reg __390301_390301;
   reg _390302_390302 ; 
   reg __390302_390302;
   reg _390303_390303 ; 
   reg __390303_390303;
   reg _390304_390304 ; 
   reg __390304_390304;
   reg _390305_390305 ; 
   reg __390305_390305;
   reg _390306_390306 ; 
   reg __390306_390306;
   reg _390307_390307 ; 
   reg __390307_390307;
   reg _390308_390308 ; 
   reg __390308_390308;
   reg _390309_390309 ; 
   reg __390309_390309;
   reg _390310_390310 ; 
   reg __390310_390310;
   reg _390311_390311 ; 
   reg __390311_390311;
   reg _390312_390312 ; 
   reg __390312_390312;
   reg _390313_390313 ; 
   reg __390313_390313;
   reg _390314_390314 ; 
   reg __390314_390314;
   reg _390315_390315 ; 
   reg __390315_390315;
   reg _390316_390316 ; 
   reg __390316_390316;
   reg _390317_390317 ; 
   reg __390317_390317;
   reg _390318_390318 ; 
   reg __390318_390318;
   reg _390319_390319 ; 
   reg __390319_390319;
   reg _390320_390320 ; 
   reg __390320_390320;
   reg _390321_390321 ; 
   reg __390321_390321;
   reg _390322_390322 ; 
   reg __390322_390322;
   reg _390323_390323 ; 
   reg __390323_390323;
   reg _390324_390324 ; 
   reg __390324_390324;
   reg _390325_390325 ; 
   reg __390325_390325;
   reg _390326_390326 ; 
   reg __390326_390326;
   reg _390327_390327 ; 
   reg __390327_390327;
   reg _390328_390328 ; 
   reg __390328_390328;
   reg _390329_390329 ; 
   reg __390329_390329;
   reg _390330_390330 ; 
   reg __390330_390330;
   reg _390331_390331 ; 
   reg __390331_390331;
   reg _390332_390332 ; 
   reg __390332_390332;
   reg _390333_390333 ; 
   reg __390333_390333;
   reg _390334_390334 ; 
   reg __390334_390334;
   reg _390335_390335 ; 
   reg __390335_390335;
   reg _390336_390336 ; 
   reg __390336_390336;
   reg _390337_390337 ; 
   reg __390337_390337;
   reg _390338_390338 ; 
   reg __390338_390338;
   reg _390339_390339 ; 
   reg __390339_390339;
   reg _390340_390340 ; 
   reg __390340_390340;
   reg _390341_390341 ; 
   reg __390341_390341;
   reg _390342_390342 ; 
   reg __390342_390342;
   reg _390343_390343 ; 
   reg __390343_390343;
   reg _390344_390344 ; 
   reg __390344_390344;
   reg _390345_390345 ; 
   reg __390345_390345;
   reg _390346_390346 ; 
   reg __390346_390346;
   reg _390347_390347 ; 
   reg __390347_390347;
   reg _390348_390348 ; 
   reg __390348_390348;
   reg _390349_390349 ; 
   reg __390349_390349;
   reg _390350_390350 ; 
   reg __390350_390350;
   reg _390351_390351 ; 
   reg __390351_390351;
   reg _390352_390352 ; 
   reg __390352_390352;
   reg _390353_390353 ; 
   reg __390353_390353;
   reg _390354_390354 ; 
   reg __390354_390354;
   reg _390355_390355 ; 
   reg __390355_390355;
   reg _390356_390356 ; 
   reg __390356_390356;
   reg _390357_390357 ; 
   reg __390357_390357;
   reg _390358_390358 ; 
   reg __390358_390358;
   reg _390359_390359 ; 
   reg __390359_390359;
   reg _390360_390360 ; 
   reg __390360_390360;
   reg _390361_390361 ; 
   reg __390361_390361;
   reg _390362_390362 ; 
   reg __390362_390362;
   reg _390363_390363 ; 
   reg __390363_390363;
   reg _390364_390364 ; 
   reg __390364_390364;
   reg _390365_390365 ; 
   reg __390365_390365;
   reg _390366_390366 ; 
   reg __390366_390366;
   reg _390367_390367 ; 
   reg __390367_390367;
   reg _390368_390368 ; 
   reg __390368_390368;
   reg _390369_390369 ; 
   reg __390369_390369;
   reg _390370_390370 ; 
   reg __390370_390370;
   reg _390371_390371 ; 
   reg __390371_390371;
   reg _390372_390372 ; 
   reg __390372_390372;
   reg _390373_390373 ; 
   reg __390373_390373;
   reg _390374_390374 ; 
   reg __390374_390374;
   reg _390375_390375 ; 
   reg __390375_390375;
   reg _390376_390376 ; 
   reg __390376_390376;
   reg _390377_390377 ; 
   reg __390377_390377;
   reg _390378_390378 ; 
   reg __390378_390378;
   reg _390379_390379 ; 
   reg __390379_390379;
   reg _390380_390380 ; 
   reg __390380_390380;
   reg _390381_390381 ; 
   reg __390381_390381;
   reg _390382_390382 ; 
   reg __390382_390382;
   reg _390383_390383 ; 
   reg __390383_390383;
   reg _390384_390384 ; 
   reg __390384_390384;
   reg _390385_390385 ; 
   reg __390385_390385;
   reg _390386_390386 ; 
   reg __390386_390386;
   reg _390387_390387 ; 
   reg __390387_390387;
   reg _390388_390388 ; 
   reg __390388_390388;
   reg _390389_390389 ; 
   reg __390389_390389;
   reg _390390_390390 ; 
   reg __390390_390390;
   reg _390391_390391 ; 
   reg __390391_390391;
   reg _390392_390392 ; 
   reg __390392_390392;
   reg _390393_390393 ; 
   reg __390393_390393;
   reg _390394_390394 ; 
   reg __390394_390394;
   reg _390395_390395 ; 
   reg __390395_390395;
   reg _390396_390396 ; 
   reg __390396_390396;
   reg _390397_390397 ; 
   reg __390397_390397;
   reg _390398_390398 ; 
   reg __390398_390398;
   reg _390399_390399 ; 
   reg __390399_390399;
   reg _390400_390400 ; 
   reg __390400_390400;
   reg _390401_390401 ; 
   reg __390401_390401;
   reg _390402_390402 ; 
   reg __390402_390402;
   reg _390403_390403 ; 
   reg __390403_390403;
   reg _390404_390404 ; 
   reg __390404_390404;
   reg _390405_390405 ; 
   reg __390405_390405;
   reg _390406_390406 ; 
   reg __390406_390406;
   reg _390407_390407 ; 
   reg __390407_390407;
   reg _390408_390408 ; 
   reg __390408_390408;
   reg _390409_390409 ; 
   reg __390409_390409;
   reg _390410_390410 ; 
   reg __390410_390410;
   reg _390411_390411 ; 
   reg __390411_390411;
   reg _390412_390412 ; 
   reg __390412_390412;
   reg _390413_390413 ; 
   reg __390413_390413;
   reg _390414_390414 ; 
   reg __390414_390414;
   reg _390415_390415 ; 
   reg __390415_390415;
   reg _390416_390416 ; 
   reg __390416_390416;
   reg _390417_390417 ; 
   reg __390417_390417;
   reg _390418_390418 ; 
   reg __390418_390418;
   reg _390419_390419 ; 
   reg __390419_390419;
   reg _390420_390420 ; 
   reg __390420_390420;
   reg _390421_390421 ; 
   reg __390421_390421;
   reg _390422_390422 ; 
   reg __390422_390422;
   reg _390423_390423 ; 
   reg __390423_390423;
   reg _390424_390424 ; 
   reg __390424_390424;
   reg _390425_390425 ; 
   reg __390425_390425;
   reg _390426_390426 ; 
   reg __390426_390426;
   reg _390427_390427 ; 
   reg __390427_390427;
   reg _390428_390428 ; 
   reg __390428_390428;
   reg _390429_390429 ; 
   reg __390429_390429;
   reg _390430_390430 ; 
   reg __390430_390430;
   reg _390431_390431 ; 
   reg __390431_390431;
   reg _390432_390432 ; 
   reg __390432_390432;
   reg _390433_390433 ; 
   reg __390433_390433;
   reg _390434_390434 ; 
   reg __390434_390434;
   reg _390435_390435 ; 
   reg __390435_390435;
   reg _390436_390436 ; 
   reg __390436_390436;
   reg _390437_390437 ; 
   reg __390437_390437;
   reg _390438_390438 ; 
   reg __390438_390438;
   reg _390439_390439 ; 
   reg __390439_390439;
   reg _390440_390440 ; 
   reg __390440_390440;
   reg _390441_390441 ; 
   reg __390441_390441;
   reg _390442_390442 ; 
   reg __390442_390442;
   reg _390443_390443 ; 
   reg __390443_390443;
   reg _390444_390444 ; 
   reg __390444_390444;
   reg _390445_390445 ; 
   reg __390445_390445;
   reg _390446_390446 ; 
   reg __390446_390446;
   reg _390447_390447 ; 
   reg __390447_390447;
   reg _390448_390448 ; 
   reg __390448_390448;
   reg _390449_390449 ; 
   reg __390449_390449;
   reg _390450_390450 ; 
   reg __390450_390450;
   reg _390451_390451 ; 
   reg __390451_390451;
   reg _390452_390452 ; 
   reg __390452_390452;
   reg _390453_390453 ; 
   reg __390453_390453;
   reg _390454_390454 ; 
   reg __390454_390454;
   reg _390455_390455 ; 
   reg __390455_390455;
   reg _390456_390456 ; 
   reg __390456_390456;
   reg _390457_390457 ; 
   reg __390457_390457;
   reg _390458_390458 ; 
   reg __390458_390458;
   reg _390459_390459 ; 
   reg __390459_390459;
   reg _390460_390460 ; 
   reg __390460_390460;
   reg _390461_390461 ; 
   reg __390461_390461;
   reg _390462_390462 ; 
   reg __390462_390462;
   reg _390463_390463 ; 
   reg __390463_390463;
   reg _390464_390464 ; 
   reg __390464_390464;
   reg _390465_390465 ; 
   reg __390465_390465;
   reg _390466_390466 ; 
   reg __390466_390466;
   reg _390467_390467 ; 
   reg __390467_390467;
   reg _390468_390468 ; 
   reg __390468_390468;
   reg _390469_390469 ; 
   reg __390469_390469;
   reg _390470_390470 ; 
   reg __390470_390470;
   reg _390471_390471 ; 
   reg __390471_390471;
   reg _390472_390472 ; 
   reg __390472_390472;
   reg _390473_390473 ; 
   reg __390473_390473;
   reg _390474_390474 ; 
   reg __390474_390474;
   reg _390475_390475 ; 
   reg __390475_390475;
   reg _390476_390476 ; 
   reg __390476_390476;
   reg _390477_390477 ; 
   reg __390477_390477;
   reg _390478_390478 ; 
   reg __390478_390478;
   reg _390479_390479 ; 
   reg __390479_390479;
   reg _390480_390480 ; 
   reg __390480_390480;
   reg _390481_390481 ; 
   reg __390481_390481;
   reg _390482_390482 ; 
   reg __390482_390482;
   reg _390483_390483 ; 
   reg __390483_390483;
   reg _390484_390484 ; 
   reg __390484_390484;
   reg _390485_390485 ; 
   reg __390485_390485;
   reg _390486_390486 ; 
   reg __390486_390486;
   reg _390487_390487 ; 
   reg __390487_390487;
   reg _390488_390488 ; 
   reg __390488_390488;
   reg _390489_390489 ; 
   reg __390489_390489;
   reg _390490_390490 ; 
   reg __390490_390490;
   reg _390491_390491 ; 
   reg __390491_390491;
   reg _390492_390492 ; 
   reg __390492_390492;
   reg _390493_390493 ; 
   reg __390493_390493;
   reg _390494_390494 ; 
   reg __390494_390494;
   reg _390495_390495 ; 
   reg __390495_390495;
   reg _390496_390496 ; 
   reg __390496_390496;
   reg _390497_390497 ; 
   reg __390497_390497;
   reg _390498_390498 ; 
   reg __390498_390498;
   reg _390499_390499 ; 
   reg __390499_390499;
   reg _390500_390500 ; 
   reg __390500_390500;
   reg _390501_390501 ; 
   reg __390501_390501;
   reg _390502_390502 ; 
   reg __390502_390502;
   reg _390503_390503 ; 
   reg __390503_390503;
   reg _390504_390504 ; 
   reg __390504_390504;
   reg _390505_390505 ; 
   reg __390505_390505;
   reg _390506_390506 ; 
   reg __390506_390506;
   reg _390507_390507 ; 
   reg __390507_390507;
   reg _390508_390508 ; 
   reg __390508_390508;
   reg _390509_390509 ; 
   reg __390509_390509;
   reg _390510_390510 ; 
   reg __390510_390510;
   reg _390511_390511 ; 
   reg __390511_390511;
   reg _390512_390512 ; 
   reg __390512_390512;
   reg _390513_390513 ; 
   reg __390513_390513;
   reg _390514_390514 ; 
   reg __390514_390514;
   reg _390515_390515 ; 
   reg __390515_390515;
   reg _390516_390516 ; 
   reg __390516_390516;
   reg _390517_390517 ; 
   reg __390517_390517;
   reg _390518_390518 ; 
   reg __390518_390518;
   reg _390519_390519 ; 
   reg __390519_390519;
   reg _390520_390520 ; 
   reg __390520_390520;
   reg _390521_390521 ; 
   reg __390521_390521;
   reg _390522_390522 ; 
   reg __390522_390522;
   reg _390523_390523 ; 
   reg __390523_390523;
   reg _390524_390524 ; 
   reg __390524_390524;
   reg _390525_390525 ; 
   reg __390525_390525;
   reg _390526_390526 ; 
   reg __390526_390526;
   reg _390527_390527 ; 
   reg __390527_390527;
   reg _390528_390528 ; 
   reg __390528_390528;
   reg _390529_390529 ; 
   reg __390529_390529;
   reg _390530_390530 ; 
   reg __390530_390530;
   reg _390531_390531 ; 
   reg __390531_390531;
   reg _390532_390532 ; 
   reg __390532_390532;
   reg _390533_390533 ; 
   reg __390533_390533;
   reg _390534_390534 ; 
   reg __390534_390534;
   reg _390535_390535 ; 
   reg __390535_390535;
   reg _390536_390536 ; 
   reg __390536_390536;
   reg _390537_390537 ; 
   reg __390537_390537;
   reg _390538_390538 ; 
   reg __390538_390538;
   reg _390539_390539 ; 
   reg __390539_390539;
   reg _390540_390540 ; 
   reg __390540_390540;
   reg _390541_390541 ; 
   reg __390541_390541;
   reg _390542_390542 ; 
   reg __390542_390542;
   reg _390543_390543 ; 
   reg __390543_390543;
   reg _390544_390544 ; 
   reg __390544_390544;
   reg _390545_390545 ; 
   reg __390545_390545;
   reg _390546_390546 ; 
   reg __390546_390546;
   reg _390547_390547 ; 
   reg __390547_390547;
   reg _390548_390548 ; 
   reg __390548_390548;
   reg _390549_390549 ; 
   reg __390549_390549;
   reg _390550_390550 ; 
   reg __390550_390550;
   reg _390551_390551 ; 
   reg __390551_390551;
   reg _390552_390552 ; 
   reg __390552_390552;
   reg _390553_390553 ; 
   reg __390553_390553;
   reg _390554_390554 ; 
   reg __390554_390554;
   reg _390555_390555 ; 
   reg __390555_390555;
   reg _390556_390556 ; 
   reg __390556_390556;
   reg _390557_390557 ; 
   reg __390557_390557;
   reg _390558_390558 ; 
   reg __390558_390558;
   reg _390559_390559 ; 
   reg __390559_390559;
   reg _390560_390560 ; 
   reg __390560_390560;
   reg _390561_390561 ; 
   reg __390561_390561;
   reg _390562_390562 ; 
   reg __390562_390562;
   reg _390563_390563 ; 
   reg __390563_390563;
   reg _390564_390564 ; 
   reg __390564_390564;
   reg _390565_390565 ; 
   reg __390565_390565;
   reg _390566_390566 ; 
   reg __390566_390566;
   reg _390567_390567 ; 
   reg __390567_390567;
   reg _390568_390568 ; 
   reg __390568_390568;
   reg _390569_390569 ; 
   reg __390569_390569;
   reg _390570_390570 ; 
   reg __390570_390570;
   reg _390571_390571 ; 
   reg __390571_390571;
   reg _390572_390572 ; 
   reg __390572_390572;
   reg _390573_390573 ; 
   reg __390573_390573;
   reg _390574_390574 ; 
   reg __390574_390574;
   reg _390575_390575 ; 
   reg __390575_390575;
   reg _390576_390576 ; 
   reg __390576_390576;
   reg _390577_390577 ; 
   reg __390577_390577;
   reg _390578_390578 ; 
   reg __390578_390578;
   reg _390579_390579 ; 
   reg __390579_390579;
   reg _390580_390580 ; 
   reg __390580_390580;
   reg _390581_390581 ; 
   reg __390581_390581;
   reg _390582_390582 ; 
   reg __390582_390582;
   reg _390583_390583 ; 
   reg __390583_390583;
   reg _390584_390584 ; 
   reg __390584_390584;
   reg _390585_390585 ; 
   reg __390585_390585;
   reg _390586_390586 ; 
   reg __390586_390586;
   reg _390587_390587 ; 
   reg __390587_390587;
   reg _390588_390588 ; 
   reg __390588_390588;
   reg _390589_390589 ; 
   reg __390589_390589;
   reg _390590_390590 ; 
   reg __390590_390590;
   reg _390591_390591 ; 
   reg __390591_390591;
   reg _390592_390592 ; 
   reg __390592_390592;
   reg _390593_390593 ; 
   reg __390593_390593;
   reg _390594_390594 ; 
   reg __390594_390594;
   reg _390595_390595 ; 
   reg __390595_390595;
   reg _390596_390596 ; 
   reg __390596_390596;
   reg _390597_390597 ; 
   reg __390597_390597;
   reg _390598_390598 ; 
   reg __390598_390598;
   reg _390599_390599 ; 
   reg __390599_390599;
   reg _390600_390600 ; 
   reg __390600_390600;
   reg _390601_390601 ; 
   reg __390601_390601;
   reg _390602_390602 ; 
   reg __390602_390602;
   reg _390603_390603 ; 
   reg __390603_390603;
   reg _390604_390604 ; 
   reg __390604_390604;
   reg _390605_390605 ; 
   reg __390605_390605;
   reg _390606_390606 ; 
   reg __390606_390606;
   reg _390607_390607 ; 
   reg __390607_390607;
   reg _390608_390608 ; 
   reg __390608_390608;
   reg _390609_390609 ; 
   reg __390609_390609;
   reg _390610_390610 ; 
   reg __390610_390610;
   reg _390611_390611 ; 
   reg __390611_390611;
   reg _390612_390612 ; 
   reg __390612_390612;
   reg _390613_390613 ; 
   reg __390613_390613;
   reg _390614_390614 ; 
   reg __390614_390614;
   reg _390615_390615 ; 
   reg __390615_390615;
   reg _390616_390616 ; 
   reg __390616_390616;
   reg _390617_390617 ; 
   reg __390617_390617;
   reg _390618_390618 ; 
   reg __390618_390618;
   reg _390619_390619 ; 
   reg __390619_390619;
   reg _390620_390620 ; 
   reg __390620_390620;
   reg _390621_390621 ; 
   reg __390621_390621;
   reg _390622_390622 ; 
   reg __390622_390622;
   reg _390623_390623 ; 
   reg __390623_390623;
   reg _390624_390624 ; 
   reg __390624_390624;
   reg _390625_390625 ; 
   reg __390625_390625;
   reg _390626_390626 ; 
   reg __390626_390626;
   reg _390627_390627 ; 
   reg __390627_390627;
   reg _390628_390628 ; 
   reg __390628_390628;
   reg _390629_390629 ; 
   reg __390629_390629;
   reg _390630_390630 ; 
   reg __390630_390630;
   reg _390631_390631 ; 
   reg __390631_390631;
   reg _390632_390632 ; 
   reg __390632_390632;
   reg _390633_390633 ; 
   reg __390633_390633;
   reg _390634_390634 ; 
   reg __390634_390634;
   reg _390635_390635 ; 
   reg __390635_390635;
   reg _390636_390636 ; 
   reg __390636_390636;
   reg _390637_390637 ; 
   reg __390637_390637;
   reg _390638_390638 ; 
   reg __390638_390638;
   reg _390639_390639 ; 
   reg __390639_390639;
   reg _390640_390640 ; 
   reg __390640_390640;
   reg _390641_390641 ; 
   reg __390641_390641;
   reg _390642_390642 ; 
   reg __390642_390642;
   reg _390643_390643 ; 
   reg __390643_390643;
   reg _390644_390644 ; 
   reg __390644_390644;
   reg _390645_390645 ; 
   reg __390645_390645;
   reg _390646_390646 ; 
   reg __390646_390646;
   reg _390647_390647 ; 
   reg __390647_390647;
   reg _390648_390648 ; 
   reg __390648_390648;
   reg _390649_390649 ; 
   reg __390649_390649;
   reg _390650_390650 ; 
   reg __390650_390650;
   reg _390651_390651 ; 
   reg __390651_390651;
   reg _390652_390652 ; 
   reg __390652_390652;
   reg _390653_390653 ; 
   reg __390653_390653;
   reg _390654_390654 ; 
   reg __390654_390654;
   reg _390655_390655 ; 
   reg __390655_390655;
   reg _390656_390656 ; 
   reg __390656_390656;
   reg _390657_390657 ; 
   reg __390657_390657;
   reg _390658_390658 ; 
   reg __390658_390658;
   reg _390659_390659 ; 
   reg __390659_390659;
   reg _390660_390660 ; 
   reg __390660_390660;
   reg _390661_390661 ; 
   reg __390661_390661;
   reg _390662_390662 ; 
   reg __390662_390662;
   reg _390663_390663 ; 
   reg __390663_390663;
   reg _390664_390664 ; 
   reg __390664_390664;
   reg _390665_390665 ; 
   reg __390665_390665;
   reg _390666_390666 ; 
   reg __390666_390666;
   reg _390667_390667 ; 
   reg __390667_390667;
   reg _390668_390668 ; 
   reg __390668_390668;
   reg _390669_390669 ; 
   reg __390669_390669;
   reg _390670_390670 ; 
   reg __390670_390670;
   reg _390671_390671 ; 
   reg __390671_390671;
   reg _390672_390672 ; 
   reg __390672_390672;
   reg _390673_390673 ; 
   reg __390673_390673;
   reg _390674_390674 ; 
   reg __390674_390674;
   reg _390675_390675 ; 
   reg __390675_390675;
   reg _390676_390676 ; 
   reg __390676_390676;
   reg _390677_390677 ; 
   reg __390677_390677;
   reg _390678_390678 ; 
   reg __390678_390678;
   reg _390679_390679 ; 
   reg __390679_390679;
   reg _390680_390680 ; 
   reg __390680_390680;
   reg _390681_390681 ; 
   reg __390681_390681;
   reg _390682_390682 ; 
   reg __390682_390682;
   reg _390683_390683 ; 
   reg __390683_390683;
   reg _390684_390684 ; 
   reg __390684_390684;
   reg _390685_390685 ; 
   reg __390685_390685;
   reg _390686_390686 ; 
   reg __390686_390686;
   reg _390687_390687 ; 
   reg __390687_390687;
   reg _390688_390688 ; 
   reg __390688_390688;
   reg _390689_390689 ; 
   reg __390689_390689;
   reg _390690_390690 ; 
   reg __390690_390690;
   reg _390691_390691 ; 
   reg __390691_390691;
   reg _390692_390692 ; 
   reg __390692_390692;
   reg _390693_390693 ; 
   reg __390693_390693;
   reg _390694_390694 ; 
   reg __390694_390694;
   reg _390695_390695 ; 
   reg __390695_390695;
   reg _390696_390696 ; 
   reg __390696_390696;
   reg _390697_390697 ; 
   reg __390697_390697;
   reg _390698_390698 ; 
   reg __390698_390698;
   reg _390699_390699 ; 
   reg __390699_390699;
   reg _390700_390700 ; 
   reg __390700_390700;
   reg _390701_390701 ; 
   reg __390701_390701;
   reg _390702_390702 ; 
   reg __390702_390702;
   reg _390703_390703 ; 
   reg __390703_390703;
   reg _390704_390704 ; 
   reg __390704_390704;
   reg _390705_390705 ; 
   reg __390705_390705;
   reg _390706_390706 ; 
   reg __390706_390706;
   reg _390707_390707 ; 
   reg __390707_390707;
   reg _390708_390708 ; 
   reg __390708_390708;
   reg _390709_390709 ; 
   reg __390709_390709;
   reg _390710_390710 ; 
   reg __390710_390710;
   reg _390711_390711 ; 
   reg __390711_390711;
   reg _390712_390712 ; 
   reg __390712_390712;
   reg _390713_390713 ; 
   reg __390713_390713;
   reg _390714_390714 ; 
   reg __390714_390714;
   reg _390715_390715 ; 
   reg __390715_390715;
   reg _390716_390716 ; 
   reg __390716_390716;
   reg _390717_390717 ; 
   reg __390717_390717;
   reg _390718_390718 ; 
   reg __390718_390718;
   reg _390719_390719 ; 
   reg __390719_390719;
   reg _390720_390720 ; 
   reg __390720_390720;
   reg _390721_390721 ; 
   reg __390721_390721;
   reg _390722_390722 ; 
   reg __390722_390722;
   reg _390723_390723 ; 
   reg __390723_390723;
   reg _390724_390724 ; 
   reg __390724_390724;
   reg _390725_390725 ; 
   reg __390725_390725;
   reg _390726_390726 ; 
   reg __390726_390726;
   reg _390727_390727 ; 
   reg __390727_390727;
   reg _390728_390728 ; 
   reg __390728_390728;
   reg _390729_390729 ; 
   reg __390729_390729;
   reg _390730_390730 ; 
   reg __390730_390730;
   reg _390731_390731 ; 
   reg __390731_390731;
   reg _390732_390732 ; 
   reg __390732_390732;
   reg _390733_390733 ; 
   reg __390733_390733;
   reg _390734_390734 ; 
   reg __390734_390734;
   reg _390735_390735 ; 
   reg __390735_390735;
   reg _390736_390736 ; 
   reg __390736_390736;
   reg _390737_390737 ; 
   reg __390737_390737;
   reg _390738_390738 ; 
   reg __390738_390738;
   reg _390739_390739 ; 
   reg __390739_390739;
   reg _390740_390740 ; 
   reg __390740_390740;
   reg _390741_390741 ; 
   reg __390741_390741;
   reg _390742_390742 ; 
   reg __390742_390742;
   reg _390743_390743 ; 
   reg __390743_390743;
   reg _390744_390744 ; 
   reg __390744_390744;
   reg _390745_390745 ; 
   reg __390745_390745;
   reg _390746_390746 ; 
   reg __390746_390746;
   reg _390747_390747 ; 
   reg __390747_390747;
   reg _390748_390748 ; 
   reg __390748_390748;
   reg _390749_390749 ; 
   reg __390749_390749;
   reg _390750_390750 ; 
   reg __390750_390750;
   reg _390751_390751 ; 
   reg __390751_390751;
   reg _390752_390752 ; 
   reg __390752_390752;
   reg _390753_390753 ; 
   reg __390753_390753;
   reg _390754_390754 ; 
   reg __390754_390754;
   reg _390755_390755 ; 
   reg __390755_390755;
   reg _390756_390756 ; 
   reg __390756_390756;
   reg _390757_390757 ; 
   reg __390757_390757;
   reg _390758_390758 ; 
   reg __390758_390758;
   reg _390759_390759 ; 
   reg __390759_390759;
   reg _390760_390760 ; 
   reg __390760_390760;
   reg _390761_390761 ; 
   reg __390761_390761;
   reg _390762_390762 ; 
   reg __390762_390762;
   reg _390763_390763 ; 
   reg __390763_390763;
   reg _390764_390764 ; 
   reg __390764_390764;
   reg _390765_390765 ; 
   reg __390765_390765;
   reg _390766_390766 ; 
   reg __390766_390766;
   reg _390767_390767 ; 
   reg __390767_390767;
   reg _390768_390768 ; 
   reg __390768_390768;
   reg _390769_390769 ; 
   reg __390769_390769;
   reg _390770_390770 ; 
   reg __390770_390770;
   reg _390771_390771 ; 
   reg __390771_390771;
   reg _390772_390772 ; 
   reg __390772_390772;
   reg _390773_390773 ; 
   reg __390773_390773;
   reg _390774_390774 ; 
   reg __390774_390774;
   reg _390775_390775 ; 
   reg __390775_390775;
   reg _390776_390776 ; 
   reg __390776_390776;
   reg _390777_390777 ; 
   reg __390777_390777;
   reg _390778_390778 ; 
   reg __390778_390778;
   reg _390779_390779 ; 
   reg __390779_390779;
   reg _390780_390780 ; 
   reg __390780_390780;
   reg _390781_390781 ; 
   reg __390781_390781;
   reg _390782_390782 ; 
   reg __390782_390782;
   reg _390783_390783 ; 
   reg __390783_390783;
   reg _390784_390784 ; 
   reg __390784_390784;
   reg _390785_390785 ; 
   reg __390785_390785;
   reg _390786_390786 ; 
   reg __390786_390786;
   reg _390787_390787 ; 
   reg __390787_390787;
   reg _390788_390788 ; 
   reg __390788_390788;
   reg _390789_390789 ; 
   reg __390789_390789;
   reg _390790_390790 ; 
   reg __390790_390790;
   reg _390791_390791 ; 
   reg __390791_390791;
   reg _390792_390792 ; 
   reg __390792_390792;
   reg _390793_390793 ; 
   reg __390793_390793;
   reg _390794_390794 ; 
   reg __390794_390794;
   reg _390795_390795 ; 
   reg __390795_390795;
   reg _390796_390796 ; 
   reg __390796_390796;
   reg _390797_390797 ; 
   reg __390797_390797;
   reg _390798_390798 ; 
   reg __390798_390798;
   reg _390799_390799 ; 
   reg __390799_390799;
   reg _390800_390800 ; 
   reg __390800_390800;
   reg _390801_390801 ; 
   reg __390801_390801;
   reg _390802_390802 ; 
   reg __390802_390802;
   reg _390803_390803 ; 
   reg __390803_390803;
   reg _390804_390804 ; 
   reg __390804_390804;
   reg _390805_390805 ; 
   reg __390805_390805;
   reg _390806_390806 ; 
   reg __390806_390806;
   reg _390807_390807 ; 
   reg __390807_390807;
   reg _390808_390808 ; 
   reg __390808_390808;
   reg _390809_390809 ; 
   reg __390809_390809;
   reg _390810_390810 ; 
   reg __390810_390810;
   reg _390811_390811 ; 
   reg __390811_390811;
   reg _390812_390812 ; 
   reg __390812_390812;
   reg _390813_390813 ; 
   reg __390813_390813;
   reg _390814_390814 ; 
   reg __390814_390814;
   reg _390815_390815 ; 
   reg __390815_390815;
   reg _390816_390816 ; 
   reg __390816_390816;
   reg _390817_390817 ; 
   reg __390817_390817;
   reg _390818_390818 ; 
   reg __390818_390818;
   reg _390819_390819 ; 
   reg __390819_390819;
   reg _390820_390820 ; 
   reg __390820_390820;
   reg _390821_390821 ; 
   reg __390821_390821;
   reg _390822_390822 ; 
   reg __390822_390822;
   reg _390823_390823 ; 
   reg __390823_390823;
   reg _390824_390824 ; 
   reg __390824_390824;
   reg _390825_390825 ; 
   reg __390825_390825;
   reg _390826_390826 ; 
   reg __390826_390826;
   reg _390827_390827 ; 
   reg __390827_390827;
   reg _390828_390828 ; 
   reg __390828_390828;
   reg _390829_390829 ; 
   reg __390829_390829;
   reg _390830_390830 ; 
   reg __390830_390830;
   reg _390831_390831 ; 
   reg __390831_390831;
   reg _390832_390832 ; 
   reg __390832_390832;
   reg _390833_390833 ; 
   reg __390833_390833;
   reg _390834_390834 ; 
   reg __390834_390834;
   reg _390835_390835 ; 
   reg __390835_390835;
   reg _390836_390836 ; 
   reg __390836_390836;
   reg _390837_390837 ; 
   reg __390837_390837;
   reg _390838_390838 ; 
   reg __390838_390838;
   reg _390839_390839 ; 
   reg __390839_390839;
   reg _390840_390840 ; 
   reg __390840_390840;
   reg _390841_390841 ; 
   reg __390841_390841;
   reg _390842_390842 ; 
   reg __390842_390842;
   reg _390843_390843 ; 
   reg __390843_390843;
   reg _390844_390844 ; 
   reg __390844_390844;
   reg _390845_390845 ; 
   reg __390845_390845;
   reg _390846_390846 ; 
   reg __390846_390846;
   reg _390847_390847 ; 
   reg __390847_390847;
   reg _390848_390848 ; 
   reg __390848_390848;
   reg _390849_390849 ; 
   reg __390849_390849;
   reg _390850_390850 ; 
   reg __390850_390850;
   reg _390851_390851 ; 
   reg __390851_390851;
   reg _390852_390852 ; 
   reg __390852_390852;
   reg _390853_390853 ; 
   reg __390853_390853;
   reg _390854_390854 ; 
   reg __390854_390854;
   reg _390855_390855 ; 
   reg __390855_390855;
   reg _390856_390856 ; 
   reg __390856_390856;
   reg _390857_390857 ; 
   reg __390857_390857;
   reg _390858_390858 ; 
   reg __390858_390858;
   reg _390859_390859 ; 
   reg __390859_390859;
   reg _390860_390860 ; 
   reg __390860_390860;
   reg _390861_390861 ; 
   reg __390861_390861;
   reg _390862_390862 ; 
   reg __390862_390862;
   reg _390863_390863 ; 
   reg __390863_390863;
   reg _390864_390864 ; 
   reg __390864_390864;
   reg _390865_390865 ; 
   reg __390865_390865;
   reg _390866_390866 ; 
   reg __390866_390866;
   reg _390867_390867 ; 
   reg __390867_390867;
   reg _390868_390868 ; 
   reg __390868_390868;
   reg _390869_390869 ; 
   reg __390869_390869;
   reg _390870_390870 ; 
   reg __390870_390870;
   reg _390871_390871 ; 
   reg __390871_390871;
   reg _390872_390872 ; 
   reg __390872_390872;
   reg _390873_390873 ; 
   reg __390873_390873;
   reg _390874_390874 ; 
   reg __390874_390874;
   reg _390875_390875 ; 
   reg __390875_390875;
   reg _390876_390876 ; 
   reg __390876_390876;
   reg _390877_390877 ; 
   reg __390877_390877;
   reg _390878_390878 ; 
   reg __390878_390878;
   reg _390879_390879 ; 
   reg __390879_390879;
   reg _390880_390880 ; 
   reg __390880_390880;
   reg _390881_390881 ; 
   reg __390881_390881;
   reg _390882_390882 ; 
   reg __390882_390882;
   reg _390883_390883 ; 
   reg __390883_390883;
   reg _390884_390884 ; 
   reg __390884_390884;
   reg _390885_390885 ; 
   reg __390885_390885;
   reg _390886_390886 ; 
   reg __390886_390886;
   reg _390887_390887 ; 
   reg __390887_390887;
   reg _390888_390888 ; 
   reg __390888_390888;
   reg _390889_390889 ; 
   reg __390889_390889;
   reg _390890_390890 ; 
   reg __390890_390890;
   reg _390891_390891 ; 
   reg __390891_390891;
   reg _390892_390892 ; 
   reg __390892_390892;
   reg _390893_390893 ; 
   reg __390893_390893;
   reg _390894_390894 ; 
   reg __390894_390894;
   reg _390895_390895 ; 
   reg __390895_390895;
   reg _390896_390896 ; 
   reg __390896_390896;
   reg _390897_390897 ; 
   reg __390897_390897;
   reg _390898_390898 ; 
   reg __390898_390898;
   reg _390899_390899 ; 
   reg __390899_390899;
   reg _390900_390900 ; 
   reg __390900_390900;
   reg _390901_390901 ; 
   reg __390901_390901;
   reg _390902_390902 ; 
   reg __390902_390902;
   reg _390903_390903 ; 
   reg __390903_390903;
   reg _390904_390904 ; 
   reg __390904_390904;
   reg _390905_390905 ; 
   reg __390905_390905;
   reg _390906_390906 ; 
   reg __390906_390906;
   reg _390907_390907 ; 
   reg __390907_390907;
   reg _390908_390908 ; 
   reg __390908_390908;
   reg _390909_390909 ; 
   reg __390909_390909;
   reg _390910_390910 ; 
   reg __390910_390910;
   reg _390911_390911 ; 
   reg __390911_390911;
   reg _390912_390912 ; 
   reg __390912_390912;
   reg _390913_390913 ; 
   reg __390913_390913;
   reg _390914_390914 ; 
   reg __390914_390914;
   reg _390915_390915 ; 
   reg __390915_390915;
   reg _390916_390916 ; 
   reg __390916_390916;
   reg _390917_390917 ; 
   reg __390917_390917;
   reg _390918_390918 ; 
   reg __390918_390918;
   reg _390919_390919 ; 
   reg __390919_390919;
   reg _390920_390920 ; 
   reg __390920_390920;
   reg _390921_390921 ; 
   reg __390921_390921;
   reg _390922_390922 ; 
   reg __390922_390922;
   reg _390923_390923 ; 
   reg __390923_390923;
   reg _390924_390924 ; 
   reg __390924_390924;
   reg _390925_390925 ; 
   reg __390925_390925;
   reg _390926_390926 ; 
   reg __390926_390926;
   reg _390927_390927 ; 
   reg __390927_390927;
   reg _390928_390928 ; 
   reg __390928_390928;
   reg _390929_390929 ; 
   reg __390929_390929;
   reg _390930_390930 ; 
   reg __390930_390930;
   reg _390931_390931 ; 
   reg __390931_390931;
   reg _390932_390932 ; 
   reg __390932_390932;
   reg _390933_390933 ; 
   reg __390933_390933;
   reg _390934_390934 ; 
   reg __390934_390934;
   reg _390935_390935 ; 
   reg __390935_390935;
   reg _390936_390936 ; 
   reg __390936_390936;
   reg _390937_390937 ; 
   reg __390937_390937;
   reg _390938_390938 ; 
   reg __390938_390938;
   reg _390939_390939 ; 
   reg __390939_390939;
   reg _390940_390940 ; 
   reg __390940_390940;
   reg _390941_390941 ; 
   reg __390941_390941;
   reg _390942_390942 ; 
   reg __390942_390942;
   reg _390943_390943 ; 
   reg __390943_390943;
   reg _390944_390944 ; 
   reg __390944_390944;
   reg _390945_390945 ; 
   reg __390945_390945;
   reg _390946_390946 ; 
   reg __390946_390946;
   reg _390947_390947 ; 
   reg __390947_390947;
   reg _390948_390948 ; 
   reg __390948_390948;
   reg _390949_390949 ; 
   reg __390949_390949;
   reg _390950_390950 ; 
   reg __390950_390950;
   reg _390951_390951 ; 
   reg __390951_390951;
   reg _390952_390952 ; 
   reg __390952_390952;
   reg _390953_390953 ; 
   reg __390953_390953;
   reg _390954_390954 ; 
   reg __390954_390954;
   reg _390955_390955 ; 
   reg __390955_390955;
   reg _390956_390956 ; 
   reg __390956_390956;
   reg _390957_390957 ; 
   reg __390957_390957;
   reg _390958_390958 ; 
   reg __390958_390958;
   reg _390959_390959 ; 
   reg __390959_390959;
   reg _390960_390960 ; 
   reg __390960_390960;
   reg _390961_390961 ; 
   reg __390961_390961;
   reg _390962_390962 ; 
   reg __390962_390962;
   reg _390963_390963 ; 
   reg __390963_390963;
   reg _390964_390964 ; 
   reg __390964_390964;
   reg _390965_390965 ; 
   reg __390965_390965;
   reg _390966_390966 ; 
   reg __390966_390966;
   reg _390967_390967 ; 
   reg __390967_390967;
   reg _390968_390968 ; 
   reg __390968_390968;
   reg _390969_390969 ; 
   reg __390969_390969;
   reg _390970_390970 ; 
   reg __390970_390970;
   reg _390971_390971 ; 
   reg __390971_390971;
   reg _390972_390972 ; 
   reg __390972_390972;
   reg _390973_390973 ; 
   reg __390973_390973;
   reg _390974_390974 ; 
   reg __390974_390974;
   reg _390975_390975 ; 
   reg __390975_390975;
   reg _390976_390976 ; 
   reg __390976_390976;
   reg _390977_390977 ; 
   reg __390977_390977;
   reg _390978_390978 ; 
   reg __390978_390978;
   reg _390979_390979 ; 
   reg __390979_390979;
   reg _390980_390980 ; 
   reg __390980_390980;
   reg _390981_390981 ; 
   reg __390981_390981;
   reg _390982_390982 ; 
   reg __390982_390982;
   reg _390983_390983 ; 
   reg __390983_390983;
   reg _390984_390984 ; 
   reg __390984_390984;
   reg _390985_390985 ; 
   reg __390985_390985;
   reg _390986_390986 ; 
   reg __390986_390986;
   reg _390987_390987 ; 
   reg __390987_390987;
   reg _390988_390988 ; 
   reg __390988_390988;
   reg _390989_390989 ; 
   reg __390989_390989;
   reg _390990_390990 ; 
   reg __390990_390990;
   reg _390991_390991 ; 
   reg __390991_390991;
   reg _390992_390992 ; 
   reg __390992_390992;
   reg _390993_390993 ; 
   reg __390993_390993;
   reg _390994_390994 ; 
   reg __390994_390994;
   reg _390995_390995 ; 
   reg __390995_390995;
   reg _390996_390996 ; 
   reg __390996_390996;
   reg _390997_390997 ; 
   reg __390997_390997;
   reg _390998_390998 ; 
   reg __390998_390998;
   reg _390999_390999 ; 
   reg __390999_390999;
   reg _391000_391000 ; 
   reg __391000_391000;
   reg _391001_391001 ; 
   reg __391001_391001;
   reg _391002_391002 ; 
   reg __391002_391002;
   reg _391003_391003 ; 
   reg __391003_391003;
   reg _391004_391004 ; 
   reg __391004_391004;
   reg _391005_391005 ; 
   reg __391005_391005;
   reg _391006_391006 ; 
   reg __391006_391006;
   reg _391007_391007 ; 
   reg __391007_391007;
   reg _391008_391008 ; 
   reg __391008_391008;
   reg _391009_391009 ; 
   reg __391009_391009;
   reg _391010_391010 ; 
   reg __391010_391010;
   reg _391011_391011 ; 
   reg __391011_391011;
   reg _391012_391012 ; 
   reg __391012_391012;
   reg _391013_391013 ; 
   reg __391013_391013;
   reg _391014_391014 ; 
   reg __391014_391014;
   reg _391015_391015 ; 
   reg __391015_391015;
   reg _391016_391016 ; 
   reg __391016_391016;
   reg _391017_391017 ; 
   reg __391017_391017;
   reg _391018_391018 ; 
   reg __391018_391018;
   reg _391019_391019 ; 
   reg __391019_391019;
   reg _391020_391020 ; 
   reg __391020_391020;
   reg _391021_391021 ; 
   reg __391021_391021;
   reg _391022_391022 ; 
   reg __391022_391022;
   reg _391023_391023 ; 
   reg __391023_391023;
   reg _391024_391024 ; 
   reg __391024_391024;
   reg _391025_391025 ; 
   reg __391025_391025;
   reg _391026_391026 ; 
   reg __391026_391026;
   reg _391027_391027 ; 
   reg __391027_391027;
   reg _391028_391028 ; 
   reg __391028_391028;
   reg _391029_391029 ; 
   reg __391029_391029;
   reg _391030_391030 ; 
   reg __391030_391030;
   reg _391031_391031 ; 
   reg __391031_391031;
   reg _391032_391032 ; 
   reg __391032_391032;
   reg _391033_391033 ; 
   reg __391033_391033;
   reg _391034_391034 ; 
   reg __391034_391034;
   reg _391035_391035 ; 
   reg __391035_391035;
   reg _391036_391036 ; 
   reg __391036_391036;
   reg _391037_391037 ; 
   reg __391037_391037;
   reg _391038_391038 ; 
   reg __391038_391038;
   reg _391039_391039 ; 
   reg __391039_391039;
   reg _391040_391040 ; 
   reg __391040_391040;
   reg _391041_391041 ; 
   reg __391041_391041;
   reg _391042_391042 ; 
   reg __391042_391042;
   reg _391043_391043 ; 
   reg __391043_391043;
   reg _391044_391044 ; 
   reg __391044_391044;
   reg _391045_391045 ; 
   reg __391045_391045;
   reg _391046_391046 ; 
   reg __391046_391046;
   reg _391047_391047 ; 
   reg __391047_391047;
   reg _391048_391048 ; 
   reg __391048_391048;
   reg _391049_391049 ; 
   reg __391049_391049;
   reg _391050_391050 ; 
   reg __391050_391050;
   reg _391051_391051 ; 
   reg __391051_391051;
   reg _391052_391052 ; 
   reg __391052_391052;
   reg _391053_391053 ; 
   reg __391053_391053;
   reg _391054_391054 ; 
   reg __391054_391054;
   reg _391055_391055 ; 
   reg __391055_391055;
   reg _391056_391056 ; 
   reg __391056_391056;
   reg _391057_391057 ; 
   reg __391057_391057;
   reg _391058_391058 ; 
   reg __391058_391058;
   reg _391059_391059 ; 
   reg __391059_391059;
   reg _391060_391060 ; 
   reg __391060_391060;
   reg _391061_391061 ; 
   reg __391061_391061;
   reg _391062_391062 ; 
   reg __391062_391062;
   reg _391063_391063 ; 
   reg __391063_391063;
   reg _391064_391064 ; 
   reg __391064_391064;
   reg _391065_391065 ; 
   reg __391065_391065;
   reg _391066_391066 ; 
   reg __391066_391066;
   reg _391067_391067 ; 
   reg __391067_391067;
   reg _391068_391068 ; 
   reg __391068_391068;
   reg _391069_391069 ; 
   reg __391069_391069;
   reg _391070_391070 ; 
   reg __391070_391070;
   reg _391071_391071 ; 
   reg __391071_391071;
   reg _391072_391072 ; 
   reg __391072_391072;
   reg _391073_391073 ; 
   reg __391073_391073;
   reg _391074_391074 ; 
   reg __391074_391074;
   reg _391075_391075 ; 
   reg __391075_391075;
   reg _391076_391076 ; 
   reg __391076_391076;
   reg _391077_391077 ; 
   reg __391077_391077;
   reg _391078_391078 ; 
   reg __391078_391078;
   reg _391079_391079 ; 
   reg __391079_391079;
   reg _391080_391080 ; 
   reg __391080_391080;
   reg _391081_391081 ; 
   reg __391081_391081;
   reg _391082_391082 ; 
   reg __391082_391082;
   reg _391083_391083 ; 
   reg __391083_391083;
   reg _391084_391084 ; 
   reg __391084_391084;
   reg _391085_391085 ; 
   reg __391085_391085;
   reg _391086_391086 ; 
   reg __391086_391086;
   reg _391087_391087 ; 
   reg __391087_391087;
   reg _391088_391088 ; 
   reg __391088_391088;
   reg _391089_391089 ; 
   reg __391089_391089;
   reg _391090_391090 ; 
   reg __391090_391090;
   reg _391091_391091 ; 
   reg __391091_391091;
   reg _391092_391092 ; 
   reg __391092_391092;
   reg _391093_391093 ; 
   reg __391093_391093;
   reg _391094_391094 ; 
   reg __391094_391094;
   reg _391095_391095 ; 
   reg __391095_391095;
   reg _391096_391096 ; 
   reg __391096_391096;
   reg _391097_391097 ; 
   reg __391097_391097;
   reg _391098_391098 ; 
   reg __391098_391098;
   reg _391099_391099 ; 
   reg __391099_391099;
   reg _391100_391100 ; 
   reg __391100_391100;
   reg _391101_391101 ; 
   reg __391101_391101;
   reg _391102_391102 ; 
   reg __391102_391102;
   reg _391103_391103 ; 
   reg __391103_391103;
   reg _391104_391104 ; 
   reg __391104_391104;
   reg _391105_391105 ; 
   reg __391105_391105;
   reg _391106_391106 ; 
   reg __391106_391106;
   reg _391107_391107 ; 
   reg __391107_391107;
   reg _391108_391108 ; 
   reg __391108_391108;
   reg _391109_391109 ; 
   reg __391109_391109;
   reg _391110_391110 ; 
   reg __391110_391110;
   reg _391111_391111 ; 
   reg __391111_391111;
   reg _391112_391112 ; 
   reg __391112_391112;
   reg _391113_391113 ; 
   reg __391113_391113;
   reg _391114_391114 ; 
   reg __391114_391114;
   reg _391115_391115 ; 
   reg __391115_391115;
   reg _391116_391116 ; 
   reg __391116_391116;
   reg _391117_391117 ; 
   reg __391117_391117;
   reg _391118_391118 ; 
   reg __391118_391118;
   reg _391119_391119 ; 
   reg __391119_391119;
   reg _391120_391120 ; 
   reg __391120_391120;
   reg _391121_391121 ; 
   reg __391121_391121;
   reg _391122_391122 ; 
   reg __391122_391122;
   reg _391123_391123 ; 
   reg __391123_391123;
   reg _391124_391124 ; 
   reg __391124_391124;
   reg _391125_391125 ; 
   reg __391125_391125;
   reg _391126_391126 ; 
   reg __391126_391126;
   reg _391127_391127 ; 
   reg __391127_391127;
   reg _391128_391128 ; 
   reg __391128_391128;
   reg _391129_391129 ; 
   reg __391129_391129;
   reg _391130_391130 ; 
   reg __391130_391130;
   reg _391131_391131 ; 
   reg __391131_391131;
   reg _391132_391132 ; 
   reg __391132_391132;
   reg _391133_391133 ; 
   reg __391133_391133;
   reg _391134_391134 ; 
   reg __391134_391134;
   reg _391135_391135 ; 
   reg __391135_391135;
   reg _391136_391136 ; 
   reg __391136_391136;
   reg _391137_391137 ; 
   reg __391137_391137;
   reg _391138_391138 ; 
   reg __391138_391138;
   reg _391139_391139 ; 
   reg __391139_391139;
   reg _391140_391140 ; 
   reg __391140_391140;
   reg _391141_391141 ; 
   reg __391141_391141;
   reg _391142_391142 ; 
   reg __391142_391142;
   reg _391143_391143 ; 
   reg __391143_391143;
   reg _391144_391144 ; 
   reg __391144_391144;
   reg _391145_391145 ; 
   reg __391145_391145;
   reg _391146_391146 ; 
   reg __391146_391146;
   reg _391147_391147 ; 
   reg __391147_391147;
   reg _391148_391148 ; 
   reg __391148_391148;
   reg _391149_391149 ; 
   reg __391149_391149;
   reg _391150_391150 ; 
   reg __391150_391150;
   reg _391151_391151 ; 
   reg __391151_391151;
   reg _391152_391152 ; 
   reg __391152_391152;
   reg _391153_391153 ; 
   reg __391153_391153;
   reg _391154_391154 ; 
   reg __391154_391154;
   reg _391155_391155 ; 
   reg __391155_391155;
   reg _391156_391156 ; 
   reg __391156_391156;
   reg _391157_391157 ; 
   reg __391157_391157;
   reg _391158_391158 ; 
   reg __391158_391158;
   reg _391159_391159 ; 
   reg __391159_391159;
   reg _391160_391160 ; 
   reg __391160_391160;
   reg _391161_391161 ; 
   reg __391161_391161;
   reg _391162_391162 ; 
   reg __391162_391162;
   reg _391163_391163 ; 
   reg __391163_391163;
   reg _391164_391164 ; 
   reg __391164_391164;
   reg _391165_391165 ; 
   reg __391165_391165;
   reg _391166_391166 ; 
   reg __391166_391166;
   reg _391167_391167 ; 
   reg __391167_391167;
   reg _391168_391168 ; 
   reg __391168_391168;
   reg _391169_391169 ; 
   reg __391169_391169;
   reg _391170_391170 ; 
   reg __391170_391170;
   reg _391171_391171 ; 
   reg __391171_391171;
   reg _391172_391172 ; 
   reg __391172_391172;
   reg _391173_391173 ; 
   reg __391173_391173;
   reg _391174_391174 ; 
   reg __391174_391174;
   reg _391175_391175 ; 
   reg __391175_391175;
   reg _391176_391176 ; 
   reg __391176_391176;
   reg _391177_391177 ; 
   reg __391177_391177;
   reg _391178_391178 ; 
   reg __391178_391178;
   reg _391179_391179 ; 
   reg __391179_391179;
   reg _391180_391180 ; 
   reg __391180_391180;
   reg _391181_391181 ; 
   reg __391181_391181;
   reg _391182_391182 ; 
   reg __391182_391182;
   reg _391183_391183 ; 
   reg __391183_391183;
   reg _391184_391184 ; 
   reg __391184_391184;
   reg _391185_391185 ; 
   reg __391185_391185;
   reg _391186_391186 ; 
   reg __391186_391186;
   reg _391187_391187 ; 
   reg __391187_391187;
   reg _391188_391188 ; 
   reg __391188_391188;
   reg _391189_391189 ; 
   reg __391189_391189;
   reg _391190_391190 ; 
   reg __391190_391190;
   reg _391191_391191 ; 
   reg __391191_391191;
   reg _391192_391192 ; 
   reg __391192_391192;
   reg _391193_391193 ; 
   reg __391193_391193;
   reg _391194_391194 ; 
   reg __391194_391194;
   reg _391195_391195 ; 
   reg __391195_391195;
   reg _391196_391196 ; 
   reg __391196_391196;
   reg _391197_391197 ; 
   reg __391197_391197;
   reg _391198_391198 ; 
   reg __391198_391198;
   reg _391199_391199 ; 
   reg __391199_391199;
   reg _391200_391200 ; 
   reg __391200_391200;
   reg _391201_391201 ; 
   reg __391201_391201;
   reg _391202_391202 ; 
   reg __391202_391202;
   reg _391203_391203 ; 
   reg __391203_391203;
   reg _391204_391204 ; 
   reg __391204_391204;
   reg _391205_391205 ; 
   reg __391205_391205;
   reg _391206_391206 ; 
   reg __391206_391206;
   reg _391207_391207 ; 
   reg __391207_391207;
   reg _391208_391208 ; 
   reg __391208_391208;
   reg _391209_391209 ; 
   reg __391209_391209;
   reg _391210_391210 ; 
   reg __391210_391210;
   reg _391211_391211 ; 
   reg __391211_391211;
   reg _391212_391212 ; 
   reg __391212_391212;
   reg _391213_391213 ; 
   reg __391213_391213;
   reg _391214_391214 ; 
   reg __391214_391214;
   reg _391215_391215 ; 
   reg __391215_391215;
   reg _391216_391216 ; 
   reg __391216_391216;
   reg _391217_391217 ; 
   reg __391217_391217;
   reg _391218_391218 ; 
   reg __391218_391218;
   reg _391219_391219 ; 
   reg __391219_391219;
   reg _391220_391220 ; 
   reg __391220_391220;
   reg _391221_391221 ; 
   reg __391221_391221;
   reg _391222_391222 ; 
   reg __391222_391222;
   reg _391223_391223 ; 
   reg __391223_391223;
   reg _391224_391224 ; 
   reg __391224_391224;
   reg _391225_391225 ; 
   reg __391225_391225;
   reg _391226_391226 ; 
   reg __391226_391226;
   reg _391227_391227 ; 
   reg __391227_391227;
   reg _391228_391228 ; 
   reg __391228_391228;
   reg _391229_391229 ; 
   reg __391229_391229;
   reg _391230_391230 ; 
   reg __391230_391230;
   reg _391231_391231 ; 
   reg __391231_391231;
   reg _391232_391232 ; 
   reg __391232_391232;
   reg _391233_391233 ; 
   reg __391233_391233;
   reg _391234_391234 ; 
   reg __391234_391234;
   reg _391235_391235 ; 
   reg __391235_391235;
   reg _391236_391236 ; 
   reg __391236_391236;
   reg _391237_391237 ; 
   reg __391237_391237;
   reg _391238_391238 ; 
   reg __391238_391238;
   reg _391239_391239 ; 
   reg __391239_391239;
   reg _391240_391240 ; 
   reg __391240_391240;
   reg _391241_391241 ; 
   reg __391241_391241;
   reg _391242_391242 ; 
   reg __391242_391242;
   reg _391243_391243 ; 
   reg __391243_391243;
   reg _391244_391244 ; 
   reg __391244_391244;
   reg _391245_391245 ; 
   reg __391245_391245;
   reg _391246_391246 ; 
   reg __391246_391246;
   reg _391247_391247 ; 
   reg __391247_391247;
   reg _391248_391248 ; 
   reg __391248_391248;
   reg _391249_391249 ; 
   reg __391249_391249;
   reg _391250_391250 ; 
   reg __391250_391250;
   reg _391251_391251 ; 
   reg __391251_391251;
   reg _391252_391252 ; 
   reg __391252_391252;
   reg _391253_391253 ; 
   reg __391253_391253;
   reg _391254_391254 ; 
   reg __391254_391254;
   reg _391255_391255 ; 
   reg __391255_391255;
   reg _391256_391256 ; 
   reg __391256_391256;
   reg _391257_391257 ; 
   reg __391257_391257;
   reg _391258_391258 ; 
   reg __391258_391258;
   reg _391259_391259 ; 
   reg __391259_391259;
   reg _391260_391260 ; 
   reg __391260_391260;
   reg _391261_391261 ; 
   reg __391261_391261;
   reg _391262_391262 ; 
   reg __391262_391262;
   reg _391263_391263 ; 
   reg __391263_391263;
   reg _391264_391264 ; 
   reg __391264_391264;
   reg _391265_391265 ; 
   reg __391265_391265;
   reg _391266_391266 ; 
   reg __391266_391266;
   reg _391267_391267 ; 
   reg __391267_391267;
   reg _391268_391268 ; 
   reg __391268_391268;
   reg _391269_391269 ; 
   reg __391269_391269;
   reg _391270_391270 ; 
   reg __391270_391270;
   reg _391271_391271 ; 
   reg __391271_391271;
   reg _391272_391272 ; 
   reg __391272_391272;
   reg _391273_391273 ; 
   reg __391273_391273;
   reg _391274_391274 ; 
   reg __391274_391274;
   reg _391275_391275 ; 
   reg __391275_391275;
   reg _391276_391276 ; 
   reg __391276_391276;
   reg _391277_391277 ; 
   reg __391277_391277;
   reg _391278_391278 ; 
   reg __391278_391278;
   reg _391279_391279 ; 
   reg __391279_391279;
   reg _391280_391280 ; 
   reg __391280_391280;
   reg _391281_391281 ; 
   reg __391281_391281;
   reg _391282_391282 ; 
   reg __391282_391282;
   reg _391283_391283 ; 
   reg __391283_391283;
   reg _391284_391284 ; 
   reg __391284_391284;
   reg _391285_391285 ; 
   reg __391285_391285;
   reg _391286_391286 ; 
   reg __391286_391286;
   reg _391287_391287 ; 
   reg __391287_391287;
   reg _391288_391288 ; 
   reg __391288_391288;
   reg _391289_391289 ; 
   reg __391289_391289;
   reg _391290_391290 ; 
   reg __391290_391290;
   reg _391291_391291 ; 
   reg __391291_391291;
   reg _391292_391292 ; 
   reg __391292_391292;
   reg _391293_391293 ; 
   reg __391293_391293;
   reg _391294_391294 ; 
   reg __391294_391294;
   reg _391295_391295 ; 
   reg __391295_391295;
   reg _391296_391296 ; 
   reg __391296_391296;
   reg _391297_391297 ; 
   reg __391297_391297;
   reg _391298_391298 ; 
   reg __391298_391298;
   reg _391299_391299 ; 
   reg __391299_391299;
   reg _391300_391300 ; 
   reg __391300_391300;
   reg _391301_391301 ; 
   reg __391301_391301;
   reg _391302_391302 ; 
   reg __391302_391302;
   reg _391303_391303 ; 
   reg __391303_391303;
   reg _391304_391304 ; 
   reg __391304_391304;
   reg _391305_391305 ; 
   reg __391305_391305;
   reg _391306_391306 ; 
   reg __391306_391306;
   reg _391307_391307 ; 
   reg __391307_391307;
   reg _391308_391308 ; 
   reg __391308_391308;
   reg _391309_391309 ; 
   reg __391309_391309;
   reg _391310_391310 ; 
   reg __391310_391310;
   reg _391311_391311 ; 
   reg __391311_391311;
   reg _391312_391312 ; 
   reg __391312_391312;
   reg _391313_391313 ; 
   reg __391313_391313;
   reg _391314_391314 ; 
   reg __391314_391314;
   reg _391315_391315 ; 
   reg __391315_391315;
   reg _391316_391316 ; 
   reg __391316_391316;
   reg _391317_391317 ; 
   reg __391317_391317;
   reg _391318_391318 ; 
   reg __391318_391318;
   reg _391319_391319 ; 
   reg __391319_391319;
   reg _391320_391320 ; 
   reg __391320_391320;
   reg _391321_391321 ; 
   reg __391321_391321;
   reg _391322_391322 ; 
   reg __391322_391322;
   reg _391323_391323 ; 
   reg __391323_391323;
   reg _391324_391324 ; 
   reg __391324_391324;
   reg _391325_391325 ; 
   reg __391325_391325;
   reg _391326_391326 ; 
   reg __391326_391326;
   reg _391327_391327 ; 
   reg __391327_391327;
   reg _391328_391328 ; 
   reg __391328_391328;
   reg _391329_391329 ; 
   reg __391329_391329;
   reg _391330_391330 ; 
   reg __391330_391330;
   reg _391331_391331 ; 
   reg __391331_391331;
   reg _391332_391332 ; 
   reg __391332_391332;
   reg _391333_391333 ; 
   reg __391333_391333;
   reg _391334_391334 ; 
   reg __391334_391334;
   reg _391335_391335 ; 
   reg __391335_391335;
   reg _391336_391336 ; 
   reg __391336_391336;
   reg _391337_391337 ; 
   reg __391337_391337;
   reg _391338_391338 ; 
   reg __391338_391338;
   reg _391339_391339 ; 
   reg __391339_391339;
   reg _391340_391340 ; 
   reg __391340_391340;
   reg _391341_391341 ; 
   reg __391341_391341;
   reg _391342_391342 ; 
   reg __391342_391342;
   reg _391343_391343 ; 
   reg __391343_391343;
   reg _391344_391344 ; 
   reg __391344_391344;
   reg _391345_391345 ; 
   reg __391345_391345;
   reg _391346_391346 ; 
   reg __391346_391346;
   reg _391347_391347 ; 
   reg __391347_391347;
   reg _391348_391348 ; 
   reg __391348_391348;
   reg _391349_391349 ; 
   reg __391349_391349;
   reg _391350_391350 ; 
   reg __391350_391350;
   reg _391351_391351 ; 
   reg __391351_391351;
   reg _391352_391352 ; 
   reg __391352_391352;
   reg _391353_391353 ; 
   reg __391353_391353;
   reg _391354_391354 ; 
   reg __391354_391354;
   reg _391355_391355 ; 
   reg __391355_391355;
   reg _391356_391356 ; 
   reg __391356_391356;
   reg _391357_391357 ; 
   reg __391357_391357;
   reg _391358_391358 ; 
   reg __391358_391358;
   reg _391359_391359 ; 
   reg __391359_391359;
   reg _391360_391360 ; 
   reg __391360_391360;
   reg _391361_391361 ; 
   reg __391361_391361;
   reg _391362_391362 ; 
   reg __391362_391362;
   reg _391363_391363 ; 
   reg __391363_391363;
   reg _391364_391364 ; 
   reg __391364_391364;
   reg _391365_391365 ; 
   reg __391365_391365;
   reg _391366_391366 ; 
   reg __391366_391366;
   reg _391367_391367 ; 
   reg __391367_391367;
   reg _391368_391368 ; 
   reg __391368_391368;
   reg _391369_391369 ; 
   reg __391369_391369;
   reg _391370_391370 ; 
   reg __391370_391370;
   reg _391371_391371 ; 
   reg __391371_391371;
   reg _391372_391372 ; 
   reg __391372_391372;
   reg _391373_391373 ; 
   reg __391373_391373;
   reg _391374_391374 ; 
   reg __391374_391374;
   reg _391375_391375 ; 
   reg __391375_391375;
   reg _391376_391376 ; 
   reg __391376_391376;
   reg _391377_391377 ; 
   reg __391377_391377;
   reg _391378_391378 ; 
   reg __391378_391378;
   reg _391379_391379 ; 
   reg __391379_391379;
   reg _391380_391380 ; 
   reg __391380_391380;
   reg _391381_391381 ; 
   reg __391381_391381;
   reg _391382_391382 ; 
   reg __391382_391382;
   reg _391383_391383 ; 
   reg __391383_391383;
   reg _391384_391384 ; 
   reg __391384_391384;
   reg _391385_391385 ; 
   reg __391385_391385;
   reg _391386_391386 ; 
   reg __391386_391386;
   reg _391387_391387 ; 
   reg __391387_391387;
   reg _391388_391388 ; 
   reg __391388_391388;
   reg _391389_391389 ; 
   reg __391389_391389;
   reg _391390_391390 ; 
   reg __391390_391390;
   reg _391391_391391 ; 
   reg __391391_391391;
   reg _391392_391392 ; 
   reg __391392_391392;
   reg _391393_391393 ; 
   reg __391393_391393;
   reg _391394_391394 ; 
   reg __391394_391394;
   reg _391395_391395 ; 
   reg __391395_391395;
   reg _391396_391396 ; 
   reg __391396_391396;
   reg _391397_391397 ; 
   reg __391397_391397;
   reg _391398_391398 ; 
   reg __391398_391398;
   reg _391399_391399 ; 
   reg __391399_391399;
   reg _391400_391400 ; 
   reg __391400_391400;
   reg _391401_391401 ; 
   reg __391401_391401;
   reg _391402_391402 ; 
   reg __391402_391402;
   reg _391403_391403 ; 
   reg __391403_391403;
   reg _391404_391404 ; 
   reg __391404_391404;
   reg _391405_391405 ; 
   reg __391405_391405;
   reg _391406_391406 ; 
   reg __391406_391406;
   reg _391407_391407 ; 
   reg __391407_391407;
   reg _391408_391408 ; 
   reg __391408_391408;
   reg _391409_391409 ; 
   reg __391409_391409;
   reg _391410_391410 ; 
   reg __391410_391410;
   reg _391411_391411 ; 
   reg __391411_391411;
   reg _391412_391412 ; 
   reg __391412_391412;
   reg _391413_391413 ; 
   reg __391413_391413;
   reg _391414_391414 ; 
   reg __391414_391414;
   reg _391415_391415 ; 
   reg __391415_391415;
   reg _391416_391416 ; 
   reg __391416_391416;
   reg _391417_391417 ; 
   reg __391417_391417;
   reg _391418_391418 ; 
   reg __391418_391418;
   reg _391419_391419 ; 
   reg __391419_391419;
   reg _391420_391420 ; 
   reg __391420_391420;
   reg _391421_391421 ; 
   reg __391421_391421;
   reg _391422_391422 ; 
   reg __391422_391422;
   reg _391423_391423 ; 
   reg __391423_391423;
   reg _391424_391424 ; 
   reg __391424_391424;
   reg _391425_391425 ; 
   reg __391425_391425;
   reg _391426_391426 ; 
   reg __391426_391426;
   reg _391427_391427 ; 
   reg __391427_391427;
   reg _391428_391428 ; 
   reg __391428_391428;
   reg _391429_391429 ; 
   reg __391429_391429;
   reg _391430_391430 ; 
   reg __391430_391430;
   reg _391431_391431 ; 
   reg __391431_391431;
   reg _391432_391432 ; 
   reg __391432_391432;
   reg _391433_391433 ; 
   reg __391433_391433;
   reg _391434_391434 ; 
   reg __391434_391434;
   reg _391435_391435 ; 
   reg __391435_391435;
   reg _391436_391436 ; 
   reg __391436_391436;
   reg _391437_391437 ; 
   reg __391437_391437;
   reg _391438_391438 ; 
   reg __391438_391438;
   reg _391439_391439 ; 
   reg __391439_391439;
   reg _391440_391440 ; 
   reg __391440_391440;
   reg _391441_391441 ; 
   reg __391441_391441;
   reg _391442_391442 ; 
   reg __391442_391442;
   reg _391443_391443 ; 
   reg __391443_391443;
   reg _391444_391444 ; 
   reg __391444_391444;
   reg _391445_391445 ; 
   reg __391445_391445;
   reg _391446_391446 ; 
   reg __391446_391446;
   reg _391447_391447 ; 
   reg __391447_391447;
   reg _391448_391448 ; 
   reg __391448_391448;
   reg _391449_391449 ; 
   reg __391449_391449;
   reg _391450_391450 ; 
   reg __391450_391450;
   reg _391451_391451 ; 
   reg __391451_391451;
   reg _391452_391452 ; 
   reg __391452_391452;
   reg _391453_391453 ; 
   reg __391453_391453;
   reg _391454_391454 ; 
   reg __391454_391454;
   reg _391455_391455 ; 
   reg __391455_391455;
   reg _391456_391456 ; 
   reg __391456_391456;
   reg _391457_391457 ; 
   reg __391457_391457;
   reg _391458_391458 ; 
   reg __391458_391458;
   reg _391459_391459 ; 
   reg __391459_391459;
   reg _391460_391460 ; 
   reg __391460_391460;
   reg _391461_391461 ; 
   reg __391461_391461;
   reg _391462_391462 ; 
   reg __391462_391462;
   reg _391463_391463 ; 
   reg __391463_391463;
   reg _391464_391464 ; 
   reg __391464_391464;
   reg _391465_391465 ; 
   reg __391465_391465;
   reg _391466_391466 ; 
   reg __391466_391466;
   reg _391467_391467 ; 
   reg __391467_391467;
   reg _391468_391468 ; 
   reg __391468_391468;
   reg _391469_391469 ; 
   reg __391469_391469;
   reg _391470_391470 ; 
   reg __391470_391470;
   reg _391471_391471 ; 
   reg __391471_391471;
   reg _391472_391472 ; 
   reg __391472_391472;
   reg _391473_391473 ; 
   reg __391473_391473;
   reg _391474_391474 ; 
   reg __391474_391474;
   reg _391475_391475 ; 
   reg __391475_391475;
   reg _391476_391476 ; 
   reg __391476_391476;
   reg _391477_391477 ; 
   reg __391477_391477;
   reg _391478_391478 ; 
   reg __391478_391478;
   reg _391479_391479 ; 
   reg __391479_391479;
   reg _391480_391480 ; 
   reg __391480_391480;
   reg _391481_391481 ; 
   reg __391481_391481;
   reg _391482_391482 ; 
   reg __391482_391482;
   reg _391483_391483 ; 
   reg __391483_391483;
   reg _391484_391484 ; 
   reg __391484_391484;
   reg _391485_391485 ; 
   reg __391485_391485;
   reg _391486_391486 ; 
   reg __391486_391486;
   reg _391487_391487 ; 
   reg __391487_391487;
   reg _391488_391488 ; 
   reg __391488_391488;
   reg _391489_391489 ; 
   reg __391489_391489;
   reg _391490_391490 ; 
   reg __391490_391490;
   reg _391491_391491 ; 
   reg __391491_391491;
   reg _391492_391492 ; 
   reg __391492_391492;
   reg _391493_391493 ; 
   reg __391493_391493;
   reg _391494_391494 ; 
   reg __391494_391494;
   reg _391495_391495 ; 
   reg __391495_391495;
   reg _391496_391496 ; 
   reg __391496_391496;
   reg _391497_391497 ; 
   reg __391497_391497;
   reg _391498_391498 ; 
   reg __391498_391498;
   reg _391499_391499 ; 
   reg __391499_391499;
   reg _391500_391500 ; 
   reg __391500_391500;
   reg _391501_391501 ; 
   reg __391501_391501;
   reg _391502_391502 ; 
   reg __391502_391502;
   reg _391503_391503 ; 
   reg __391503_391503;
   reg _391504_391504 ; 
   reg __391504_391504;
   reg _391505_391505 ; 
   reg __391505_391505;
   reg _391506_391506 ; 
   reg __391506_391506;
   reg _391507_391507 ; 
   reg __391507_391507;
   reg _391508_391508 ; 
   reg __391508_391508;
   reg _391509_391509 ; 
   reg __391509_391509;
   reg _391510_391510 ; 
   reg __391510_391510;
   reg _391511_391511 ; 
   reg __391511_391511;
   reg _391512_391512 ; 
   reg __391512_391512;
   reg _391513_391513 ; 
   reg __391513_391513;
   reg _391514_391514 ; 
   reg __391514_391514;
   reg _391515_391515 ; 
   reg __391515_391515;
   reg _391516_391516 ; 
   reg __391516_391516;
   reg _391517_391517 ; 
   reg __391517_391517;
   reg _391518_391518 ; 
   reg __391518_391518;
   reg _391519_391519 ; 
   reg __391519_391519;
   reg _391520_391520 ; 
   reg __391520_391520;
   reg _391521_391521 ; 
   reg __391521_391521;
   reg _391522_391522 ; 
   reg __391522_391522;
   reg _391523_391523 ; 
   reg __391523_391523;
   reg _391524_391524 ; 
   reg __391524_391524;
   reg _391525_391525 ; 
   reg __391525_391525;
   reg _391526_391526 ; 
   reg __391526_391526;
   reg _391527_391527 ; 
   reg __391527_391527;
   reg _391528_391528 ; 
   reg __391528_391528;
   reg _391529_391529 ; 
   reg __391529_391529;
   reg _391530_391530 ; 
   reg __391530_391530;
   reg _391531_391531 ; 
   reg __391531_391531;
   reg _391532_391532 ; 
   reg __391532_391532;
   reg _391533_391533 ; 
   reg __391533_391533;
   reg _391534_391534 ; 
   reg __391534_391534;
   reg _391535_391535 ; 
   reg __391535_391535;
   reg _391536_391536 ; 
   reg __391536_391536;
   reg _391537_391537 ; 
   reg __391537_391537;
   reg _391538_391538 ; 
   reg __391538_391538;
   reg _391539_391539 ; 
   reg __391539_391539;
   reg _391540_391540 ; 
   reg __391540_391540;
   reg _391541_391541 ; 
   reg __391541_391541;
   reg _391542_391542 ; 
   reg __391542_391542;
   reg _391543_391543 ; 
   reg __391543_391543;
   reg _391544_391544 ; 
   reg __391544_391544;
   reg _391545_391545 ; 
   reg __391545_391545;
   reg _391546_391546 ; 
   reg __391546_391546;
   reg _391547_391547 ; 
   reg __391547_391547;
   reg _391548_391548 ; 
   reg __391548_391548;
   reg _391549_391549 ; 
   reg __391549_391549;
   reg _391550_391550 ; 
   reg __391550_391550;
   reg _391551_391551 ; 
   reg __391551_391551;
   reg _391552_391552 ; 
   reg __391552_391552;
   reg _391553_391553 ; 
   reg __391553_391553;
   reg _391554_391554 ; 
   reg __391554_391554;
   reg _391555_391555 ; 
   reg __391555_391555;
   reg _391556_391556 ; 
   reg __391556_391556;
   reg _391557_391557 ; 
   reg __391557_391557;
   reg _391558_391558 ; 
   reg __391558_391558;
   reg _391559_391559 ; 
   reg __391559_391559;
   reg _391560_391560 ; 
   reg __391560_391560;
   reg _391561_391561 ; 
   reg __391561_391561;
   reg _391562_391562 ; 
   reg __391562_391562;
   reg _391563_391563 ; 
   reg __391563_391563;
   reg _391564_391564 ; 
   reg __391564_391564;
   reg _391565_391565 ; 
   reg __391565_391565;
   reg _391566_391566 ; 
   reg __391566_391566;
   reg _391567_391567 ; 
   reg __391567_391567;
   reg _391568_391568 ; 
   reg __391568_391568;
   reg _391569_391569 ; 
   reg __391569_391569;
   reg _391570_391570 ; 
   reg __391570_391570;
   reg _391571_391571 ; 
   reg __391571_391571;
   reg _391572_391572 ; 
   reg __391572_391572;
   reg _391573_391573 ; 
   reg __391573_391573;
   reg _391574_391574 ; 
   reg __391574_391574;
   reg _391575_391575 ; 
   reg __391575_391575;
   reg _391576_391576 ; 
   reg __391576_391576;
   reg _391577_391577 ; 
   reg __391577_391577;
   reg _391578_391578 ; 
   reg __391578_391578;
   reg _391579_391579 ; 
   reg __391579_391579;
   reg _391580_391580 ; 
   reg __391580_391580;
   reg _391581_391581 ; 
   reg __391581_391581;
   reg _391582_391582 ; 
   reg __391582_391582;
   reg _391583_391583 ; 
   reg __391583_391583;
   reg _391584_391584 ; 
   reg __391584_391584;
   reg _391585_391585 ; 
   reg __391585_391585;
   reg _391586_391586 ; 
   reg __391586_391586;
   reg _391587_391587 ; 
   reg __391587_391587;
   reg _391588_391588 ; 
   reg __391588_391588;
   reg _391589_391589 ; 
   reg __391589_391589;
   reg _391590_391590 ; 
   reg __391590_391590;
   reg _391591_391591 ; 
   reg __391591_391591;
   reg _391592_391592 ; 
   reg __391592_391592;
   reg _391593_391593 ; 
   reg __391593_391593;
   reg _391594_391594 ; 
   reg __391594_391594;
   reg _391595_391595 ; 
   reg __391595_391595;
   reg _391596_391596 ; 
   reg __391596_391596;
   reg _391597_391597 ; 
   reg __391597_391597;
   reg _391598_391598 ; 
   reg __391598_391598;
   reg _391599_391599 ; 
   reg __391599_391599;
   reg _391600_391600 ; 
   reg __391600_391600;
   reg _391601_391601 ; 
   reg __391601_391601;
   reg _391602_391602 ; 
   reg __391602_391602;
   reg _391603_391603 ; 
   reg __391603_391603;
   reg _391604_391604 ; 
   reg __391604_391604;
   reg _391605_391605 ; 
   reg __391605_391605;
   reg _391606_391606 ; 
   reg __391606_391606;
   reg _391607_391607 ; 
   reg __391607_391607;
   reg _391608_391608 ; 
   reg __391608_391608;
   reg _391609_391609 ; 
   reg __391609_391609;
   reg _391610_391610 ; 
   reg __391610_391610;
   reg _391611_391611 ; 
   reg __391611_391611;
   reg _391612_391612 ; 
   reg __391612_391612;
   reg _391613_391613 ; 
   reg __391613_391613;
   reg _391614_391614 ; 
   reg __391614_391614;
   reg _391615_391615 ; 
   reg __391615_391615;
   reg _391616_391616 ; 
   reg __391616_391616;
   reg _391617_391617 ; 
   reg __391617_391617;
   reg _391618_391618 ; 
   reg __391618_391618;
   reg _391619_391619 ; 
   reg __391619_391619;
   reg _391620_391620 ; 
   reg __391620_391620;
   reg _391621_391621 ; 
   reg __391621_391621;
   reg _391622_391622 ; 
   reg __391622_391622;
   reg _391623_391623 ; 
   reg __391623_391623;
   reg _391624_391624 ; 
   reg __391624_391624;
   reg _391625_391625 ; 
   reg __391625_391625;
   reg _391626_391626 ; 
   reg __391626_391626;
   reg _391627_391627 ; 
   reg __391627_391627;
   reg _391628_391628 ; 
   reg __391628_391628;
   reg _391629_391629 ; 
   reg __391629_391629;
   reg _391630_391630 ; 
   reg __391630_391630;
   reg _391631_391631 ; 
   reg __391631_391631;
   reg _391632_391632 ; 
   reg __391632_391632;
   reg _391633_391633 ; 
   reg __391633_391633;
   reg _391634_391634 ; 
   reg __391634_391634;
   reg _391635_391635 ; 
   reg __391635_391635;
   reg _391636_391636 ; 
   reg __391636_391636;
   reg _391637_391637 ; 
   reg __391637_391637;
   reg _391638_391638 ; 
   reg __391638_391638;
   reg _391639_391639 ; 
   reg __391639_391639;
   reg _391640_391640 ; 
   reg __391640_391640;
   reg _391641_391641 ; 
   reg __391641_391641;
   reg _391642_391642 ; 
   reg __391642_391642;
   reg _391643_391643 ; 
   reg __391643_391643;
   reg _391644_391644 ; 
   reg __391644_391644;
   reg _391645_391645 ; 
   reg __391645_391645;
   reg _391646_391646 ; 
   reg __391646_391646;
   reg _391647_391647 ; 
   reg __391647_391647;
   reg _391648_391648 ; 
   reg __391648_391648;
   reg _391649_391649 ; 
   reg __391649_391649;
   reg _391650_391650 ; 
   reg __391650_391650;
   reg _391651_391651 ; 
   reg __391651_391651;
   reg _391652_391652 ; 
   reg __391652_391652;
   reg _391653_391653 ; 
   reg __391653_391653;
   reg _391654_391654 ; 
   reg __391654_391654;
   reg _391655_391655 ; 
   reg __391655_391655;
   reg _391656_391656 ; 
   reg __391656_391656;
   reg _391657_391657 ; 
   reg __391657_391657;
   reg _391658_391658 ; 
   reg __391658_391658;
   reg _391659_391659 ; 
   reg __391659_391659;
   reg _391660_391660 ; 
   reg __391660_391660;
   reg _391661_391661 ; 
   reg __391661_391661;
   reg _391662_391662 ; 
   reg __391662_391662;
   reg _391663_391663 ; 
   reg __391663_391663;
   reg _391664_391664 ; 
   reg __391664_391664;
   reg _391665_391665 ; 
   reg __391665_391665;
   reg _391666_391666 ; 
   reg __391666_391666;
   reg _391667_391667 ; 
   reg __391667_391667;
   reg _391668_391668 ; 
   reg __391668_391668;
   reg _391669_391669 ; 
   reg __391669_391669;
   reg _391670_391670 ; 
   reg __391670_391670;
   reg _391671_391671 ; 
   reg __391671_391671;
   reg _391672_391672 ; 
   reg __391672_391672;
   reg _391673_391673 ; 
   reg __391673_391673;
   reg _391674_391674 ; 
   reg __391674_391674;
   reg _391675_391675 ; 
   reg __391675_391675;
   reg _391676_391676 ; 
   reg __391676_391676;
   reg _391677_391677 ; 
   reg __391677_391677;
   reg _391678_391678 ; 
   reg __391678_391678;
   reg _391679_391679 ; 
   reg __391679_391679;
   reg _391680_391680 ; 
   reg __391680_391680;
   reg _391681_391681 ; 
   reg __391681_391681;
   reg _391682_391682 ; 
   reg __391682_391682;
   reg _391683_391683 ; 
   reg __391683_391683;
   reg _391684_391684 ; 
   reg __391684_391684;
   reg _391685_391685 ; 
   reg __391685_391685;
   reg _391686_391686 ; 
   reg __391686_391686;
   reg _391687_391687 ; 
   reg __391687_391687;
   reg _391688_391688 ; 
   reg __391688_391688;
   reg _391689_391689 ; 
   reg __391689_391689;
   reg _391690_391690 ; 
   reg __391690_391690;
   reg _391691_391691 ; 
   reg __391691_391691;
   reg _391692_391692 ; 
   reg __391692_391692;
   reg _391693_391693 ; 
   reg __391693_391693;
   reg _391694_391694 ; 
   reg __391694_391694;
   reg _391695_391695 ; 
   reg __391695_391695;
   reg _391696_391696 ; 
   reg __391696_391696;
   reg _391697_391697 ; 
   reg __391697_391697;
   reg _391698_391698 ; 
   reg __391698_391698;
   reg _391699_391699 ; 
   reg __391699_391699;
   reg _391700_391700 ; 
   reg __391700_391700;
   reg _391701_391701 ; 
   reg __391701_391701;
   reg _391702_391702 ; 
   reg __391702_391702;
   reg _391703_391703 ; 
   reg __391703_391703;
   reg _391704_391704 ; 
   reg __391704_391704;
   reg _391705_391705 ; 
   reg __391705_391705;
   reg _391706_391706 ; 
   reg __391706_391706;
   reg _391707_391707 ; 
   reg __391707_391707;
   reg _391708_391708 ; 
   reg __391708_391708;
   reg _391709_391709 ; 
   reg __391709_391709;
   reg _391710_391710 ; 
   reg __391710_391710;
   reg _391711_391711 ; 
   reg __391711_391711;
   reg _391712_391712 ; 
   reg __391712_391712;
   reg _391713_391713 ; 
   reg __391713_391713;
   reg _391714_391714 ; 
   reg __391714_391714;
   reg _391715_391715 ; 
   reg __391715_391715;
   reg _391716_391716 ; 
   reg __391716_391716;
   reg _391717_391717 ; 
   reg __391717_391717;
   reg _391718_391718 ; 
   reg __391718_391718;
   reg _391719_391719 ; 
   reg __391719_391719;
   reg _391720_391720 ; 
   reg __391720_391720;
   reg _391721_391721 ; 
   reg __391721_391721;
   reg _391722_391722 ; 
   reg __391722_391722;
   reg _391723_391723 ; 
   reg __391723_391723;
   reg _391724_391724 ; 
   reg __391724_391724;
   reg _391725_391725 ; 
   reg __391725_391725;
   reg _391726_391726 ; 
   reg __391726_391726;
   reg _391727_391727 ; 
   reg __391727_391727;
   reg _391728_391728 ; 
   reg __391728_391728;
   reg _391729_391729 ; 
   reg __391729_391729;
   reg _391730_391730 ; 
   reg __391730_391730;
   reg _391731_391731 ; 
   reg __391731_391731;
   reg _391732_391732 ; 
   reg __391732_391732;
   reg _391733_391733 ; 
   reg __391733_391733;
   reg _391734_391734 ; 
   reg __391734_391734;
   reg _391735_391735 ; 
   reg __391735_391735;
   reg _391736_391736 ; 
   reg __391736_391736;
   reg _391737_391737 ; 
   reg __391737_391737;
   reg _391738_391738 ; 
   reg __391738_391738;
   reg _391739_391739 ; 
   reg __391739_391739;
   reg _391740_391740 ; 
   reg __391740_391740;
   reg _391741_391741 ; 
   reg __391741_391741;
   reg _391742_391742 ; 
   reg __391742_391742;
   reg _391743_391743 ; 
   reg __391743_391743;
   reg _391744_391744 ; 
   reg __391744_391744;
   reg _391745_391745 ; 
   reg __391745_391745;
   reg _391746_391746 ; 
   reg __391746_391746;
   reg _391747_391747 ; 
   reg __391747_391747;
   reg _391748_391748 ; 
   reg __391748_391748;
   reg _391749_391749 ; 
   reg __391749_391749;
   reg _391750_391750 ; 
   reg __391750_391750;
   reg _391751_391751 ; 
   reg __391751_391751;
   reg _391752_391752 ; 
   reg __391752_391752;
   reg _391753_391753 ; 
   reg __391753_391753;
   reg _391754_391754 ; 
   reg __391754_391754;
   reg _391755_391755 ; 
   reg __391755_391755;
   reg _391756_391756 ; 
   reg __391756_391756;
   reg _391757_391757 ; 
   reg __391757_391757;
   reg _391758_391758 ; 
   reg __391758_391758;
   reg _391759_391759 ; 
   reg __391759_391759;
   reg _391760_391760 ; 
   reg __391760_391760;
   reg _391761_391761 ; 
   reg __391761_391761;
   reg _391762_391762 ; 
   reg __391762_391762;
   reg _391763_391763 ; 
   reg __391763_391763;
   reg _391764_391764 ; 
   reg __391764_391764;
   reg _391765_391765 ; 
   reg __391765_391765;
   reg _391766_391766 ; 
   reg __391766_391766;
   reg _391767_391767 ; 
   reg __391767_391767;
   reg _391768_391768 ; 
   reg __391768_391768;
   reg _391769_391769 ; 
   reg __391769_391769;
   reg _391770_391770 ; 
   reg __391770_391770;
   reg _391771_391771 ; 
   reg __391771_391771;
   reg _391772_391772 ; 
   reg __391772_391772;
   reg _391773_391773 ; 
   reg __391773_391773;
   reg _391774_391774 ; 
   reg __391774_391774;
   reg _391775_391775 ; 
   reg __391775_391775;
   reg _391776_391776 ; 
   reg __391776_391776;
   reg _391777_391777 ; 
   reg __391777_391777;
   reg _391778_391778 ; 
   reg __391778_391778;
   reg _391779_391779 ; 
   reg __391779_391779;
   reg _391780_391780 ; 
   reg __391780_391780;
   reg _391781_391781 ; 
   reg __391781_391781;
   reg _391782_391782 ; 
   reg __391782_391782;
   reg _391783_391783 ; 
   reg __391783_391783;
   reg _391784_391784 ; 
   reg __391784_391784;
   reg _391785_391785 ; 
   reg __391785_391785;
   reg _391786_391786 ; 
   reg __391786_391786;
   reg _391787_391787 ; 
   reg __391787_391787;
   reg _391788_391788 ; 
   reg __391788_391788;
   reg _391789_391789 ; 
   reg __391789_391789;
   reg _391790_391790 ; 
   reg __391790_391790;
   reg _391791_391791 ; 
   reg __391791_391791;
   reg _391792_391792 ; 
   reg __391792_391792;
   reg _391793_391793 ; 
   reg __391793_391793;
   reg _391794_391794 ; 
   reg __391794_391794;
   reg _391795_391795 ; 
   reg __391795_391795;
   reg _391796_391796 ; 
   reg __391796_391796;
   reg _391797_391797 ; 
   reg __391797_391797;
   reg _391798_391798 ; 
   reg __391798_391798;
   reg _391799_391799 ; 
   reg __391799_391799;
   reg _391800_391800 ; 
   reg __391800_391800;
   reg _391801_391801 ; 
   reg __391801_391801;
   reg _391802_391802 ; 
   reg __391802_391802;
   reg _391803_391803 ; 
   reg __391803_391803;
   reg _391804_391804 ; 
   reg __391804_391804;
   reg _391805_391805 ; 
   reg __391805_391805;
   reg _391806_391806 ; 
   reg __391806_391806;
   reg _391807_391807 ; 
   reg __391807_391807;
   reg _391808_391808 ; 
   reg __391808_391808;
   reg _391809_391809 ; 
   reg __391809_391809;
   reg _391810_391810 ; 
   reg __391810_391810;
   reg _391811_391811 ; 
   reg __391811_391811;
   reg _391812_391812 ; 
   reg __391812_391812;
   reg _391813_391813 ; 
   reg __391813_391813;
   reg _391814_391814 ; 
   reg __391814_391814;
   reg _391815_391815 ; 
   reg __391815_391815;
   reg _391816_391816 ; 
   reg __391816_391816;
   reg _391817_391817 ; 
   reg __391817_391817;
   reg _391818_391818 ; 
   reg __391818_391818;
   reg _391819_391819 ; 
   reg __391819_391819;
   reg _391820_391820 ; 
   reg __391820_391820;
   reg _391821_391821 ; 
   reg __391821_391821;
   reg _391822_391822 ; 
   reg __391822_391822;
   reg _391823_391823 ; 
   reg __391823_391823;
   reg _391824_391824 ; 
   reg __391824_391824;
   reg _391825_391825 ; 
   reg __391825_391825;
   reg _391826_391826 ; 
   reg __391826_391826;
   reg _391827_391827 ; 
   reg __391827_391827;
   reg _391828_391828 ; 
   reg __391828_391828;
   reg _391829_391829 ; 
   reg __391829_391829;
   reg _391830_391830 ; 
   reg __391830_391830;
   reg _391831_391831 ; 
   reg __391831_391831;
   reg _391832_391832 ; 
   reg __391832_391832;
   reg _391833_391833 ; 
   reg __391833_391833;
   reg _391834_391834 ; 
   reg __391834_391834;
   reg _391835_391835 ; 
   reg __391835_391835;
   reg _391836_391836 ; 
   reg __391836_391836;
   reg _391837_391837 ; 
   reg __391837_391837;
   reg _391838_391838 ; 
   reg __391838_391838;
   reg _391839_391839 ; 
   reg __391839_391839;
   reg _391840_391840 ; 
   reg __391840_391840;
   reg _391841_391841 ; 
   reg __391841_391841;
   reg _391842_391842 ; 
   reg __391842_391842;
   reg _391843_391843 ; 
   reg __391843_391843;
   reg _391844_391844 ; 
   reg __391844_391844;
   reg _391845_391845 ; 
   reg __391845_391845;
   reg _391846_391846 ; 
   reg __391846_391846;
   reg _391847_391847 ; 
   reg __391847_391847;
   reg _391848_391848 ; 
   reg __391848_391848;
   reg _391849_391849 ; 
   reg __391849_391849;
   reg _391850_391850 ; 
   reg __391850_391850;
   reg _391851_391851 ; 
   reg __391851_391851;
   reg _391852_391852 ; 
   reg __391852_391852;
   reg _391853_391853 ; 
   reg __391853_391853;
   reg _391854_391854 ; 
   reg __391854_391854;
   reg _391855_391855 ; 
   reg __391855_391855;
   reg _391856_391856 ; 
   reg __391856_391856;
   reg _391857_391857 ; 
   reg __391857_391857;
   reg _391858_391858 ; 
   reg __391858_391858;
   reg _391859_391859 ; 
   reg __391859_391859;
   reg _391860_391860 ; 
   reg __391860_391860;
   reg _391861_391861 ; 
   reg __391861_391861;
   reg _391862_391862 ; 
   reg __391862_391862;
   reg _391863_391863 ; 
   reg __391863_391863;
   reg _391864_391864 ; 
   reg __391864_391864;
   reg _391865_391865 ; 
   reg __391865_391865;
   reg _391866_391866 ; 
   reg __391866_391866;
   reg _391867_391867 ; 
   reg __391867_391867;
   reg _391868_391868 ; 
   reg __391868_391868;
   reg _391869_391869 ; 
   reg __391869_391869;
   reg _391870_391870 ; 
   reg __391870_391870;
   reg _391871_391871 ; 
   reg __391871_391871;
   reg _391872_391872 ; 
   reg __391872_391872;
   reg _391873_391873 ; 
   reg __391873_391873;
   reg _391874_391874 ; 
   reg __391874_391874;
   reg _391875_391875 ; 
   reg __391875_391875;
   reg _391876_391876 ; 
   reg __391876_391876;
   reg _391877_391877 ; 
   reg __391877_391877;
   reg _391878_391878 ; 
   reg __391878_391878;
   reg _391879_391879 ; 
   reg __391879_391879;
   reg _391880_391880 ; 
   reg __391880_391880;
   reg _391881_391881 ; 
   reg __391881_391881;
   reg _391882_391882 ; 
   reg __391882_391882;
   reg _391883_391883 ; 
   reg __391883_391883;
   reg _391884_391884 ; 
   reg __391884_391884;
   reg _391885_391885 ; 
   reg __391885_391885;
   reg _391886_391886 ; 
   reg __391886_391886;
   reg _391887_391887 ; 
   reg __391887_391887;
   reg _391888_391888 ; 
   reg __391888_391888;
   reg _391889_391889 ; 
   reg __391889_391889;
   reg _391890_391890 ; 
   reg __391890_391890;
   reg _391891_391891 ; 
   reg __391891_391891;
   reg _391892_391892 ; 
   reg __391892_391892;
   reg _391893_391893 ; 
   reg __391893_391893;
   reg _391894_391894 ; 
   reg __391894_391894;
   reg _391895_391895 ; 
   reg __391895_391895;
   reg _391896_391896 ; 
   reg __391896_391896;
   reg _391897_391897 ; 
   reg __391897_391897;
   reg _391898_391898 ; 
   reg __391898_391898;
   reg _391899_391899 ; 
   reg __391899_391899;
   reg _391900_391900 ; 
   reg __391900_391900;
   reg _391901_391901 ; 
   reg __391901_391901;
   reg _391902_391902 ; 
   reg __391902_391902;
   reg _391903_391903 ; 
   reg __391903_391903;
   reg _391904_391904 ; 
   reg __391904_391904;
   reg _391905_391905 ; 
   reg __391905_391905;
   reg _391906_391906 ; 
   reg __391906_391906;
   reg _391907_391907 ; 
   reg __391907_391907;
   reg _391908_391908 ; 
   reg __391908_391908;
   reg _391909_391909 ; 
   reg __391909_391909;
   reg _391910_391910 ; 
   reg __391910_391910;
   reg _391911_391911 ; 
   reg __391911_391911;
   reg _391912_391912 ; 
   reg __391912_391912;
   reg _391913_391913 ; 
   reg __391913_391913;
   reg _391914_391914 ; 
   reg __391914_391914;
   reg _391915_391915 ; 
   reg __391915_391915;
   reg _391916_391916 ; 
   reg __391916_391916;
   reg _391917_391917 ; 
   reg __391917_391917;
   reg _391918_391918 ; 
   reg __391918_391918;
   reg _391919_391919 ; 
   reg __391919_391919;
   reg _391920_391920 ; 
   reg __391920_391920;
   reg _391921_391921 ; 
   reg __391921_391921;
   reg _391922_391922 ; 
   reg __391922_391922;
   reg _391923_391923 ; 
   reg __391923_391923;
   reg _391924_391924 ; 
   reg __391924_391924;
   reg _391925_391925 ; 
   reg __391925_391925;
   reg _391926_391926 ; 
   reg __391926_391926;
   reg _391927_391927 ; 
   reg __391927_391927;
   reg _391928_391928 ; 
   reg __391928_391928;
   reg _391929_391929 ; 
   reg __391929_391929;
   reg _391930_391930 ; 
   reg __391930_391930;
   reg _391931_391931 ; 
   reg __391931_391931;
   reg _391932_391932 ; 
   reg __391932_391932;
   reg _391933_391933 ; 
   reg __391933_391933;
   reg _391934_391934 ; 
   reg __391934_391934;
   reg _391935_391935 ; 
   reg __391935_391935;
   reg _391936_391936 ; 
   reg __391936_391936;
   reg _391937_391937 ; 
   reg __391937_391937;
   reg _391938_391938 ; 
   reg __391938_391938;
   reg _391939_391939 ; 
   reg __391939_391939;
   reg _391940_391940 ; 
   reg __391940_391940;
   reg _391941_391941 ; 
   reg __391941_391941;
   reg _391942_391942 ; 
   reg __391942_391942;
   reg _391943_391943 ; 
   reg __391943_391943;
   reg _391944_391944 ; 
   reg __391944_391944;
   reg _391945_391945 ; 
   reg __391945_391945;
   reg _391946_391946 ; 
   reg __391946_391946;
   reg _391947_391947 ; 
   reg __391947_391947;
   reg _391948_391948 ; 
   reg __391948_391948;
   reg _391949_391949 ; 
   reg __391949_391949;
   reg _391950_391950 ; 
   reg __391950_391950;
   reg _391951_391951 ; 
   reg __391951_391951;
   reg _391952_391952 ; 
   reg __391952_391952;
   reg _391953_391953 ; 
   reg __391953_391953;
   reg _391954_391954 ; 
   reg __391954_391954;
   reg _391955_391955 ; 
   reg __391955_391955;
   reg _391956_391956 ; 
   reg __391956_391956;
   reg _391957_391957 ; 
   reg __391957_391957;
   reg _391958_391958 ; 
   reg __391958_391958;
   reg _391959_391959 ; 
   reg __391959_391959;
   reg _391960_391960 ; 
   reg __391960_391960;
   reg _391961_391961 ; 
   reg __391961_391961;
   reg _391962_391962 ; 
   reg __391962_391962;
   reg _391963_391963 ; 
   reg __391963_391963;
   reg _391964_391964 ; 
   reg __391964_391964;
   reg _391965_391965 ; 
   reg __391965_391965;
   reg _391966_391966 ; 
   reg __391966_391966;
   reg _391967_391967 ; 
   reg __391967_391967;
   reg _391968_391968 ; 
   reg __391968_391968;
   reg _391969_391969 ; 
   reg __391969_391969;
   reg _391970_391970 ; 
   reg __391970_391970;
   reg _391971_391971 ; 
   reg __391971_391971;
   reg _391972_391972 ; 
   reg __391972_391972;
   reg _391973_391973 ; 
   reg __391973_391973;
   reg _391974_391974 ; 
   reg __391974_391974;
   reg _391975_391975 ; 
   reg __391975_391975;
   reg _391976_391976 ; 
   reg __391976_391976;
   reg _391977_391977 ; 
   reg __391977_391977;
   reg _391978_391978 ; 
   reg __391978_391978;
   reg _391979_391979 ; 
   reg __391979_391979;
   reg _391980_391980 ; 
   reg __391980_391980;
   reg _391981_391981 ; 
   reg __391981_391981;
   reg _391982_391982 ; 
   reg __391982_391982;
   reg _391983_391983 ; 
   reg __391983_391983;
   reg _391984_391984 ; 
   reg __391984_391984;
   reg _391985_391985 ; 
   reg __391985_391985;
   reg _391986_391986 ; 
   reg __391986_391986;
   reg _391987_391987 ; 
   reg __391987_391987;
   reg _391988_391988 ; 
   reg __391988_391988;
   reg _391989_391989 ; 
   reg __391989_391989;
   reg _391990_391990 ; 
   reg __391990_391990;
   reg _391991_391991 ; 
   reg __391991_391991;
   reg _391992_391992 ; 
   reg __391992_391992;
   reg _391993_391993 ; 
   reg __391993_391993;
   reg _391994_391994 ; 
   reg __391994_391994;
   reg _391995_391995 ; 
   reg __391995_391995;
   reg _391996_391996 ; 
   reg __391996_391996;
   reg _391997_391997 ; 
   reg __391997_391997;
   reg _391998_391998 ; 
   reg __391998_391998;
   reg _391999_391999 ; 
   reg __391999_391999;
   reg _392000_392000 ; 
   reg __392000_392000;
   reg _392001_392001 ; 
   reg __392001_392001;
   reg _392002_392002 ; 
   reg __392002_392002;
   reg _392003_392003 ; 
   reg __392003_392003;
   reg _392004_392004 ; 
   reg __392004_392004;
   reg _392005_392005 ; 
   reg __392005_392005;
   reg _392006_392006 ; 
   reg __392006_392006;
   reg _392007_392007 ; 
   reg __392007_392007;
   reg _392008_392008 ; 
   reg __392008_392008;
   reg _392009_392009 ; 
   reg __392009_392009;
   reg _392010_392010 ; 
   reg __392010_392010;
   reg _392011_392011 ; 
   reg __392011_392011;
   reg _392012_392012 ; 
   reg __392012_392012;
   reg _392013_392013 ; 
   reg __392013_392013;
   reg _392014_392014 ; 
   reg __392014_392014;
   reg _392015_392015 ; 
   reg __392015_392015;
   reg _392016_392016 ; 
   reg __392016_392016;
   reg _392017_392017 ; 
   reg __392017_392017;
   reg _392018_392018 ; 
   reg __392018_392018;
   reg _392019_392019 ; 
   reg __392019_392019;
   reg _392020_392020 ; 
   reg __392020_392020;
   reg _392021_392021 ; 
   reg __392021_392021;
   reg _392022_392022 ; 
   reg __392022_392022;
   reg _392023_392023 ; 
   reg __392023_392023;
   reg _392024_392024 ; 
   reg __392024_392024;
   reg _392025_392025 ; 
   reg __392025_392025;
   reg _392026_392026 ; 
   reg __392026_392026;
   reg _392027_392027 ; 
   reg __392027_392027;
   reg _392028_392028 ; 
   reg __392028_392028;
   reg _392029_392029 ; 
   reg __392029_392029;
   reg _392030_392030 ; 
   reg __392030_392030;
   reg _392031_392031 ; 
   reg __392031_392031;
   reg _392032_392032 ; 
   reg __392032_392032;
   reg _392033_392033 ; 
   reg __392033_392033;
   reg _392034_392034 ; 
   reg __392034_392034;
   reg _392035_392035 ; 
   reg __392035_392035;
   reg _392036_392036 ; 
   reg __392036_392036;
   reg _392037_392037 ; 
   reg __392037_392037;
   reg _392038_392038 ; 
   reg __392038_392038;
   reg _392039_392039 ; 
   reg __392039_392039;
   reg _392040_392040 ; 
   reg __392040_392040;
   reg _392041_392041 ; 
   reg __392041_392041;
   reg _392042_392042 ; 
   reg __392042_392042;
   reg _392043_392043 ; 
   reg __392043_392043;
   reg _392044_392044 ; 
   reg __392044_392044;
   reg _392045_392045 ; 
   reg __392045_392045;
   reg _392046_392046 ; 
   reg __392046_392046;
   reg _392047_392047 ; 
   reg __392047_392047;
   reg _392048_392048 ; 
   reg __392048_392048;
   reg _392049_392049 ; 
   reg __392049_392049;
   reg _392050_392050 ; 
   reg __392050_392050;
   reg _392051_392051 ; 
   reg __392051_392051;
   reg _392052_392052 ; 
   reg __392052_392052;
   reg _392053_392053 ; 
   reg __392053_392053;
   reg _392054_392054 ; 
   reg __392054_392054;
   reg _392055_392055 ; 
   reg __392055_392055;
   reg _392056_392056 ; 
   reg __392056_392056;
   reg _392057_392057 ; 
   reg __392057_392057;
   reg _392058_392058 ; 
   reg __392058_392058;
   reg _392059_392059 ; 
   reg __392059_392059;
   reg _392060_392060 ; 
   reg __392060_392060;
   reg _392061_392061 ; 
   reg __392061_392061;
   reg _392062_392062 ; 
   reg __392062_392062;
   reg _392063_392063 ; 
   reg __392063_392063;
   reg _392064_392064 ; 
   reg __392064_392064;
   reg _392065_392065 ; 
   reg __392065_392065;
   reg _392066_392066 ; 
   reg __392066_392066;
   reg _392067_392067 ; 
   reg __392067_392067;
   reg _392068_392068 ; 
   reg __392068_392068;
   reg _392069_392069 ; 
   reg __392069_392069;
   reg _392070_392070 ; 
   reg __392070_392070;
   reg _392071_392071 ; 
   reg __392071_392071;
   reg _392072_392072 ; 
   reg __392072_392072;
   reg _392073_392073 ; 
   reg __392073_392073;
   reg _392074_392074 ; 
   reg __392074_392074;
   reg _392075_392075 ; 
   reg __392075_392075;
   reg _392076_392076 ; 
   reg __392076_392076;
   reg _392077_392077 ; 
   reg __392077_392077;
   reg _392078_392078 ; 
   reg __392078_392078;
   reg _392079_392079 ; 
   reg __392079_392079;
   reg _392080_392080 ; 
   reg __392080_392080;
   reg _392081_392081 ; 
   reg __392081_392081;
   reg _392082_392082 ; 
   reg __392082_392082;
   reg _392083_392083 ; 
   reg __392083_392083;
   reg _392084_392084 ; 
   reg __392084_392084;
   reg _392085_392085 ; 
   reg __392085_392085;
   reg _392086_392086 ; 
   reg __392086_392086;
   reg _392087_392087 ; 
   reg __392087_392087;
   reg _392088_392088 ; 
   reg __392088_392088;
   reg _392089_392089 ; 
   reg __392089_392089;
   reg _392090_392090 ; 
   reg __392090_392090;
   reg _392091_392091 ; 
   reg __392091_392091;
   reg _392092_392092 ; 
   reg __392092_392092;
   reg _392093_392093 ; 
   reg __392093_392093;
   reg _392094_392094 ; 
   reg __392094_392094;
   reg _392095_392095 ; 
   reg __392095_392095;
   reg _392096_392096 ; 
   reg __392096_392096;
   reg _392097_392097 ; 
   reg __392097_392097;
   reg _392098_392098 ; 
   reg __392098_392098;
   reg _392099_392099 ; 
   reg __392099_392099;
   reg _392100_392100 ; 
   reg __392100_392100;
   reg _392101_392101 ; 
   reg __392101_392101;
   reg _392102_392102 ; 
   reg __392102_392102;
   reg _392103_392103 ; 
   reg __392103_392103;
   reg _392104_392104 ; 
   reg __392104_392104;
   reg _392105_392105 ; 
   reg __392105_392105;
   reg _392106_392106 ; 
   reg __392106_392106;
   reg _392107_392107 ; 
   reg __392107_392107;
   reg _392108_392108 ; 
   reg __392108_392108;
   reg _392109_392109 ; 
   reg __392109_392109;
   reg _392110_392110 ; 
   reg __392110_392110;
   reg _392111_392111 ; 
   reg __392111_392111;
   reg _392112_392112 ; 
   reg __392112_392112;
   reg _392113_392113 ; 
   reg __392113_392113;
   reg _392114_392114 ; 
   reg __392114_392114;
   reg _392115_392115 ; 
   reg __392115_392115;
   reg _392116_392116 ; 
   reg __392116_392116;
   reg _392117_392117 ; 
   reg __392117_392117;
   reg _392118_392118 ; 
   reg __392118_392118;
   reg _392119_392119 ; 
   reg __392119_392119;
   reg _392120_392120 ; 
   reg __392120_392120;
   reg _392121_392121 ; 
   reg __392121_392121;
   reg _392122_392122 ; 
   reg __392122_392122;
   reg _392123_392123 ; 
   reg __392123_392123;
   reg _392124_392124 ; 
   reg __392124_392124;
   reg _392125_392125 ; 
   reg __392125_392125;
   reg _392126_392126 ; 
   reg __392126_392126;
   reg _392127_392127 ; 
   reg __392127_392127;
   reg _392128_392128 ; 
   reg __392128_392128;
   reg _392129_392129 ; 
   reg __392129_392129;
   reg _392130_392130 ; 
   reg __392130_392130;
   reg _392131_392131 ; 
   reg __392131_392131;
   reg _392132_392132 ; 
   reg __392132_392132;
   reg _392133_392133 ; 
   reg __392133_392133;
   reg _392134_392134 ; 
   reg __392134_392134;
   reg _392135_392135 ; 
   reg __392135_392135;
   reg _392136_392136 ; 
   reg __392136_392136;
   reg _392137_392137 ; 
   reg __392137_392137;
   reg _392138_392138 ; 
   reg __392138_392138;
   reg _392139_392139 ; 
   reg __392139_392139;
   reg _392140_392140 ; 
   reg __392140_392140;
   reg _392141_392141 ; 
   reg __392141_392141;
   reg _392142_392142 ; 
   reg __392142_392142;
   reg _392143_392143 ; 
   reg __392143_392143;
   reg _392144_392144 ; 
   reg __392144_392144;
   reg _392145_392145 ; 
   reg __392145_392145;
   reg _392146_392146 ; 
   reg __392146_392146;
   reg _392147_392147 ; 
   reg __392147_392147;
   reg _392148_392148 ; 
   reg __392148_392148;
   reg _392149_392149 ; 
   reg __392149_392149;
   reg _392150_392150 ; 
   reg __392150_392150;
   reg _392151_392151 ; 
   reg __392151_392151;
   reg _392152_392152 ; 
   reg __392152_392152;
   reg _392153_392153 ; 
   reg __392153_392153;
   reg _392154_392154 ; 
   reg __392154_392154;
   reg _392155_392155 ; 
   reg __392155_392155;
   reg _392156_392156 ; 
   reg __392156_392156;
   reg _392157_392157 ; 
   reg __392157_392157;
   reg _392158_392158 ; 
   reg __392158_392158;
   reg _392159_392159 ; 
   reg __392159_392159;
   reg _392160_392160 ; 
   reg __392160_392160;
   reg _392161_392161 ; 
   reg __392161_392161;
   reg _392162_392162 ; 
   reg __392162_392162;
   reg _392163_392163 ; 
   reg __392163_392163;
   reg _392164_392164 ; 
   reg __392164_392164;
   reg _392165_392165 ; 
   reg __392165_392165;
   reg _392166_392166 ; 
   reg __392166_392166;
   reg _392167_392167 ; 
   reg __392167_392167;
   reg _392168_392168 ; 
   reg __392168_392168;
   reg _392169_392169 ; 
   reg __392169_392169;
   reg _392170_392170 ; 
   reg __392170_392170;
   reg _392171_392171 ; 
   reg __392171_392171;
   reg _392172_392172 ; 
   reg __392172_392172;
   reg _392173_392173 ; 
   reg __392173_392173;
   reg _392174_392174 ; 
   reg __392174_392174;
   reg _392175_392175 ; 
   reg __392175_392175;
   reg _392176_392176 ; 
   reg __392176_392176;
   reg _392177_392177 ; 
   reg __392177_392177;
   reg _392178_392178 ; 
   reg __392178_392178;
   reg _392179_392179 ; 
   reg __392179_392179;
   reg _392180_392180 ; 
   reg __392180_392180;
   reg _392181_392181 ; 
   reg __392181_392181;
   reg _392182_392182 ; 
   reg __392182_392182;
   reg _392183_392183 ; 
   reg __392183_392183;
   reg _392184_392184 ; 
   reg __392184_392184;
   reg _392185_392185 ; 
   reg __392185_392185;
   reg _392186_392186 ; 
   reg __392186_392186;
   reg _392187_392187 ; 
   reg __392187_392187;
   reg _392188_392188 ; 
   reg __392188_392188;
   reg _392189_392189 ; 
   reg __392189_392189;
   reg _392190_392190 ; 
   reg __392190_392190;
   reg _392191_392191 ; 
   reg __392191_392191;
   reg _392192_392192 ; 
   reg __392192_392192;
   reg _392193_392193 ; 
   reg __392193_392193;
   reg _392194_392194 ; 
   reg __392194_392194;
   reg _392195_392195 ; 
   reg __392195_392195;
   reg _392196_392196 ; 
   reg __392196_392196;
   reg _392197_392197 ; 
   reg __392197_392197;
   reg _392198_392198 ; 
   reg __392198_392198;
   reg _392199_392199 ; 
   reg __392199_392199;
   reg _392200_392200 ; 
   reg __392200_392200;
   reg _392201_392201 ; 
   reg __392201_392201;
   reg _392202_392202 ; 
   reg __392202_392202;
   reg _392203_392203 ; 
   reg __392203_392203;
   reg _392204_392204 ; 
   reg __392204_392204;
   reg _392205_392205 ; 
   reg __392205_392205;
   reg _392206_392206 ; 
   reg __392206_392206;
   reg _392207_392207 ; 
   reg __392207_392207;
   reg _392208_392208 ; 
   reg __392208_392208;
   reg _392209_392209 ; 
   reg __392209_392209;
   reg _392210_392210 ; 
   reg __392210_392210;
   reg _392211_392211 ; 
   reg __392211_392211;
   reg _392212_392212 ; 
   reg __392212_392212;
   reg _392213_392213 ; 
   reg __392213_392213;
   reg _392214_392214 ; 
   reg __392214_392214;
   reg _392215_392215 ; 
   reg __392215_392215;
   reg _392216_392216 ; 
   reg __392216_392216;
   reg _392217_392217 ; 
   reg __392217_392217;
   reg _392218_392218 ; 
   reg __392218_392218;
   reg _392219_392219 ; 
   reg __392219_392219;
   reg _392220_392220 ; 
   reg __392220_392220;
   reg _392221_392221 ; 
   reg __392221_392221;
   reg _392222_392222 ; 
   reg __392222_392222;
   reg _392223_392223 ; 
   reg __392223_392223;
   reg _392224_392224 ; 
   reg __392224_392224;
   reg _392225_392225 ; 
   reg __392225_392225;
   reg _392226_392226 ; 
   reg __392226_392226;
   reg _392227_392227 ; 
   reg __392227_392227;
   reg _392228_392228 ; 
   reg __392228_392228;
   reg _392229_392229 ; 
   reg __392229_392229;
   reg _392230_392230 ; 
   reg __392230_392230;
   reg _392231_392231 ; 
   reg __392231_392231;
   reg _392232_392232 ; 
   reg __392232_392232;
   reg _392233_392233 ; 
   reg __392233_392233;
   reg _392234_392234 ; 
   reg __392234_392234;
   reg _392235_392235 ; 
   reg __392235_392235;
   reg _392236_392236 ; 
   reg __392236_392236;
   reg _392237_392237 ; 
   reg __392237_392237;
   reg _392238_392238 ; 
   reg __392238_392238;
   reg _392239_392239 ; 
   reg __392239_392239;
   reg _392240_392240 ; 
   reg __392240_392240;
   reg _392241_392241 ; 
   reg __392241_392241;
   reg _392242_392242 ; 
   reg __392242_392242;
   reg _392243_392243 ; 
   reg __392243_392243;
   reg _392244_392244 ; 
   reg __392244_392244;
   reg _392245_392245 ; 
   reg __392245_392245;
   reg _392246_392246 ; 
   reg __392246_392246;
   reg _392247_392247 ; 
   reg __392247_392247;
   reg _392248_392248 ; 
   reg __392248_392248;
   reg _392249_392249 ; 
   reg __392249_392249;
   reg _392250_392250 ; 
   reg __392250_392250;
   reg _392251_392251 ; 
   reg __392251_392251;
   reg _392252_392252 ; 
   reg __392252_392252;
   reg _392253_392253 ; 
   reg __392253_392253;
   reg _392254_392254 ; 
   reg __392254_392254;
   reg _392255_392255 ; 
   reg __392255_392255;
   reg _392256_392256 ; 
   reg __392256_392256;
   reg _392257_392257 ; 
   reg __392257_392257;
   reg _392258_392258 ; 
   reg __392258_392258;
   reg _392259_392259 ; 
   reg __392259_392259;
   reg _392260_392260 ; 
   reg __392260_392260;
   reg _392261_392261 ; 
   reg __392261_392261;
   reg _392262_392262 ; 
   reg __392262_392262;
   reg _392263_392263 ; 
   reg __392263_392263;
   reg _392264_392264 ; 
   reg __392264_392264;
   reg _392265_392265 ; 
   reg __392265_392265;
   reg _392266_392266 ; 
   reg __392266_392266;
   reg _392267_392267 ; 
   reg __392267_392267;
   reg _392268_392268 ; 
   reg __392268_392268;
   reg _392269_392269 ; 
   reg __392269_392269;
   reg _392270_392270 ; 
   reg __392270_392270;
   reg _392271_392271 ; 
   reg __392271_392271;
   reg _392272_392272 ; 
   reg __392272_392272;
   reg _392273_392273 ; 
   reg __392273_392273;
   reg _392274_392274 ; 
   reg __392274_392274;
   reg _392275_392275 ; 
   reg __392275_392275;
   reg _392276_392276 ; 
   reg __392276_392276;
   reg _392277_392277 ; 
   reg __392277_392277;
   reg _392278_392278 ; 
   reg __392278_392278;
   reg _392279_392279 ; 
   reg __392279_392279;
   reg _392280_392280 ; 
   reg __392280_392280;
   reg _392281_392281 ; 
   reg __392281_392281;
   reg _392282_392282 ; 
   reg __392282_392282;
   reg _392283_392283 ; 
   reg __392283_392283;
   reg _392284_392284 ; 
   reg __392284_392284;
   reg _392285_392285 ; 
   reg __392285_392285;
   reg _392286_392286 ; 
   reg __392286_392286;
   reg _392287_392287 ; 
   reg __392287_392287;
   reg _392288_392288 ; 
   reg __392288_392288;
   reg _392289_392289 ; 
   reg __392289_392289;
   reg _392290_392290 ; 
   reg __392290_392290;
   reg _392291_392291 ; 
   reg __392291_392291;
   reg _392292_392292 ; 
   reg __392292_392292;
   reg _392293_392293 ; 
   reg __392293_392293;
   reg _392294_392294 ; 
   reg __392294_392294;
   reg _392295_392295 ; 
   reg __392295_392295;
   reg _392296_392296 ; 
   reg __392296_392296;
   reg _392297_392297 ; 
   reg __392297_392297;
   reg _392298_392298 ; 
   reg __392298_392298;
   reg _392299_392299 ; 
   reg __392299_392299;
   reg _392300_392300 ; 
   reg __392300_392300;
   reg _392301_392301 ; 
   reg __392301_392301;
   reg _392302_392302 ; 
   reg __392302_392302;
   reg _392303_392303 ; 
   reg __392303_392303;
   reg _392304_392304 ; 
   reg __392304_392304;
   reg _392305_392305 ; 
   reg __392305_392305;
   reg _392306_392306 ; 
   reg __392306_392306;
   reg _392307_392307 ; 
   reg __392307_392307;
   reg _392308_392308 ; 
   reg __392308_392308;
   reg _392309_392309 ; 
   reg __392309_392309;
   reg _392310_392310 ; 
   reg __392310_392310;
   reg _392311_392311 ; 
   reg __392311_392311;
   reg _392312_392312 ; 
   reg __392312_392312;
   reg _392313_392313 ; 
   reg __392313_392313;
   reg _392314_392314 ; 
   reg __392314_392314;
   reg _392315_392315 ; 
   reg __392315_392315;
   reg _392316_392316 ; 
   reg __392316_392316;
   reg _392317_392317 ; 
   reg __392317_392317;
   reg _392318_392318 ; 
   reg __392318_392318;
   reg _392319_392319 ; 
   reg __392319_392319;
   reg _392320_392320 ; 
   reg __392320_392320;
   reg _392321_392321 ; 
   reg __392321_392321;
   reg _392322_392322 ; 
   reg __392322_392322;
   reg _392323_392323 ; 
   reg __392323_392323;
   reg _392324_392324 ; 
   reg __392324_392324;
   reg _392325_392325 ; 
   reg __392325_392325;
   reg _392326_392326 ; 
   reg __392326_392326;
   reg _392327_392327 ; 
   reg __392327_392327;
   reg _392328_392328 ; 
   reg __392328_392328;
   reg _392329_392329 ; 
   reg __392329_392329;
   reg _392330_392330 ; 
   reg __392330_392330;
   reg _392331_392331 ; 
   reg __392331_392331;
   reg _392332_392332 ; 
   reg __392332_392332;
   reg _392333_392333 ; 
   reg __392333_392333;
   reg _392334_392334 ; 
   reg __392334_392334;
   reg _392335_392335 ; 
   reg __392335_392335;
   reg _392336_392336 ; 
   reg __392336_392336;
   reg _392337_392337 ; 
   reg __392337_392337;
   reg _392338_392338 ; 
   reg __392338_392338;
   reg _392339_392339 ; 
   reg __392339_392339;
   reg _392340_392340 ; 
   reg __392340_392340;
   reg _392341_392341 ; 
   reg __392341_392341;
   reg _392342_392342 ; 
   reg __392342_392342;
   reg _392343_392343 ; 
   reg __392343_392343;
   reg _392344_392344 ; 
   reg __392344_392344;
   reg _392345_392345 ; 
   reg __392345_392345;
   reg _392346_392346 ; 
   reg __392346_392346;
   reg _392347_392347 ; 
   reg __392347_392347;
   reg _392348_392348 ; 
   reg __392348_392348;
   reg _392349_392349 ; 
   reg __392349_392349;
   reg _392350_392350 ; 
   reg __392350_392350;
   reg _392351_392351 ; 
   reg __392351_392351;
   reg _392352_392352 ; 
   reg __392352_392352;
   reg _392353_392353 ; 
   reg __392353_392353;
   reg _392354_392354 ; 
   reg __392354_392354;
   reg _392355_392355 ; 
   reg __392355_392355;
   reg _392356_392356 ; 
   reg __392356_392356;
   reg _392357_392357 ; 
   reg __392357_392357;
   reg _392358_392358 ; 
   reg __392358_392358;
   reg _392359_392359 ; 
   reg __392359_392359;
   reg _392360_392360 ; 
   reg __392360_392360;
   reg _392361_392361 ; 
   reg __392361_392361;
   reg _392362_392362 ; 
   reg __392362_392362;
   reg _392363_392363 ; 
   reg __392363_392363;
   reg _392364_392364 ; 
   reg __392364_392364;
   reg _392365_392365 ; 
   reg __392365_392365;
   reg _392366_392366 ; 
   reg __392366_392366;
   reg _392367_392367 ; 
   reg __392367_392367;
   reg _392368_392368 ; 
   reg __392368_392368;
   reg _392369_392369 ; 
   reg __392369_392369;
   reg _392370_392370 ; 
   reg __392370_392370;
   reg _392371_392371 ; 
   reg __392371_392371;
   reg _392372_392372 ; 
   reg __392372_392372;
   reg _392373_392373 ; 
   reg __392373_392373;
   reg _392374_392374 ; 
   reg __392374_392374;
   reg _392375_392375 ; 
   reg __392375_392375;
   reg _392376_392376 ; 
   reg __392376_392376;
   reg _392377_392377 ; 
   reg __392377_392377;
   reg _392378_392378 ; 
   reg __392378_392378;
   reg _392379_392379 ; 
   reg __392379_392379;
   reg _392380_392380 ; 
   reg __392380_392380;
   reg _392381_392381 ; 
   reg __392381_392381;
   reg _392382_392382 ; 
   reg __392382_392382;
   reg _392383_392383 ; 
   reg __392383_392383;
   reg _392384_392384 ; 
   reg __392384_392384;
   reg _392385_392385 ; 
   reg __392385_392385;
   reg _392386_392386 ; 
   reg __392386_392386;
   reg _392387_392387 ; 
   reg __392387_392387;
   reg _392388_392388 ; 
   reg __392388_392388;
   reg _392389_392389 ; 
   reg __392389_392389;
   reg _392390_392390 ; 
   reg __392390_392390;
   reg _392391_392391 ; 
   reg __392391_392391;
   reg _392392_392392 ; 
   reg __392392_392392;
   reg _392393_392393 ; 
   reg __392393_392393;
   reg _392394_392394 ; 
   reg __392394_392394;
   reg _392395_392395 ; 
   reg __392395_392395;
   reg _392396_392396 ; 
   reg __392396_392396;
   reg _392397_392397 ; 
   reg __392397_392397;
   reg _392398_392398 ; 
   reg __392398_392398;
   reg _392399_392399 ; 
   reg __392399_392399;
   reg _392400_392400 ; 
   reg __392400_392400;
   reg _392401_392401 ; 
   reg __392401_392401;
   reg _392402_392402 ; 
   reg __392402_392402;
   reg _392403_392403 ; 
   reg __392403_392403;
   reg _392404_392404 ; 
   reg __392404_392404;
   reg _392405_392405 ; 
   reg __392405_392405;
   reg _392406_392406 ; 
   reg __392406_392406;
   reg _392407_392407 ; 
   reg __392407_392407;
   reg _392408_392408 ; 
   reg __392408_392408;
   reg _392409_392409 ; 
   reg __392409_392409;
   reg _392410_392410 ; 
   reg __392410_392410;
   reg _392411_392411 ; 
   reg __392411_392411;
   reg _392412_392412 ; 
   reg __392412_392412;
   reg _392413_392413 ; 
   reg __392413_392413;
   reg _392414_392414 ; 
   reg __392414_392414;
   reg _392415_392415 ; 
   reg __392415_392415;
   reg _392416_392416 ; 
   reg __392416_392416;
   reg _392417_392417 ; 
   reg __392417_392417;
   reg _392418_392418 ; 
   reg __392418_392418;
   reg _392419_392419 ; 
   reg __392419_392419;
   reg _392420_392420 ; 
   reg __392420_392420;
   reg _392421_392421 ; 
   reg __392421_392421;
   reg _392422_392422 ; 
   reg __392422_392422;
   reg _392423_392423 ; 
   reg __392423_392423;
   reg _392424_392424 ; 
   reg __392424_392424;
   reg _392425_392425 ; 
   reg __392425_392425;
   reg _392426_392426 ; 
   reg __392426_392426;
   reg _392427_392427 ; 
   reg __392427_392427;
   reg _392428_392428 ; 
   reg __392428_392428;
   reg _392429_392429 ; 
   reg __392429_392429;
   reg _392430_392430 ; 
   reg __392430_392430;
   reg _392431_392431 ; 
   reg __392431_392431;
   reg _392432_392432 ; 
   reg __392432_392432;
   reg _392433_392433 ; 
   reg __392433_392433;
   reg _392434_392434 ; 
   reg __392434_392434;
   reg _392435_392435 ; 
   reg __392435_392435;
   reg _392436_392436 ; 
   reg __392436_392436;
   reg _392437_392437 ; 
   reg __392437_392437;
   reg _392438_392438 ; 
   reg __392438_392438;
   reg _392439_392439 ; 
   reg __392439_392439;
   reg _392440_392440 ; 
   reg __392440_392440;
   reg _392441_392441 ; 
   reg __392441_392441;
   reg _392442_392442 ; 
   reg __392442_392442;
   reg _392443_392443 ; 
   reg __392443_392443;
   reg _392444_392444 ; 
   reg __392444_392444;
   reg _392445_392445 ; 
   reg __392445_392445;
   reg _392446_392446 ; 
   reg __392446_392446;
   reg _392447_392447 ; 
   reg __392447_392447;
   reg _392448_392448 ; 
   reg __392448_392448;
   reg _392449_392449 ; 
   reg __392449_392449;
   reg _392450_392450 ; 
   reg __392450_392450;
   reg _392451_392451 ; 
   reg __392451_392451;
   reg _392452_392452 ; 
   reg __392452_392452;
   reg _392453_392453 ; 
   reg __392453_392453;
   reg _392454_392454 ; 
   reg __392454_392454;
   reg _392455_392455 ; 
   reg __392455_392455;
   reg _392456_392456 ; 
   reg __392456_392456;
   reg _392457_392457 ; 
   reg __392457_392457;
   reg _392458_392458 ; 
   reg __392458_392458;
   reg _392459_392459 ; 
   reg __392459_392459;
   reg _392460_392460 ; 
   reg __392460_392460;
   reg _392461_392461 ; 
   reg __392461_392461;
   reg _392462_392462 ; 
   reg __392462_392462;
   reg _392463_392463 ; 
   reg __392463_392463;
   reg _392464_392464 ; 
   reg __392464_392464;
   reg _392465_392465 ; 
   reg __392465_392465;
   reg _392466_392466 ; 
   reg __392466_392466;
   reg _392467_392467 ; 
   reg __392467_392467;
   reg _392468_392468 ; 
   reg __392468_392468;
   reg _392469_392469 ; 
   reg __392469_392469;
   reg _392470_392470 ; 
   reg __392470_392470;
   reg _392471_392471 ; 
   reg __392471_392471;
   reg _392472_392472 ; 
   reg __392472_392472;
   reg _392473_392473 ; 
   reg __392473_392473;
   reg _392474_392474 ; 
   reg __392474_392474;
   reg _392475_392475 ; 
   reg __392475_392475;
   reg _392476_392476 ; 
   reg __392476_392476;
   reg _392477_392477 ; 
   reg __392477_392477;
   reg _392478_392478 ; 
   reg __392478_392478;
   reg _392479_392479 ; 
   reg __392479_392479;
   reg _392480_392480 ; 
   reg __392480_392480;
   reg _392481_392481 ; 
   reg __392481_392481;
   reg _392482_392482 ; 
   reg __392482_392482;
   reg _392483_392483 ; 
   reg __392483_392483;
   reg _392484_392484 ; 
   reg __392484_392484;
   reg _392485_392485 ; 
   reg __392485_392485;
   reg _392486_392486 ; 
   reg __392486_392486;
   reg _392487_392487 ; 
   reg __392487_392487;
   reg _392488_392488 ; 
   reg __392488_392488;
   reg _392489_392489 ; 
   reg __392489_392489;
   reg _392490_392490 ; 
   reg __392490_392490;
   reg _392491_392491 ; 
   reg __392491_392491;
   reg _392492_392492 ; 
   reg __392492_392492;
   reg _392493_392493 ; 
   reg __392493_392493;
   reg _392494_392494 ; 
   reg __392494_392494;
   reg _392495_392495 ; 
   reg __392495_392495;
   reg _392496_392496 ; 
   reg __392496_392496;
   reg _392497_392497 ; 
   reg __392497_392497;
   reg _392498_392498 ; 
   reg __392498_392498;
   reg _392499_392499 ; 
   reg __392499_392499;
   reg _392500_392500 ; 
   reg __392500_392500;
   reg _392501_392501 ; 
   reg __392501_392501;
   reg _392502_392502 ; 
   reg __392502_392502;
   reg _392503_392503 ; 
   reg __392503_392503;
   reg _392504_392504 ; 
   reg __392504_392504;
   reg _392505_392505 ; 
   reg __392505_392505;
   reg _392506_392506 ; 
   reg __392506_392506;
   reg _392507_392507 ; 
   reg __392507_392507;
   reg _392508_392508 ; 
   reg __392508_392508;
   reg _392509_392509 ; 
   reg __392509_392509;
   reg _392510_392510 ; 
   reg __392510_392510;
   reg _392511_392511 ; 
   reg __392511_392511;
   reg _392512_392512 ; 
   reg __392512_392512;
   reg _392513_392513 ; 
   reg __392513_392513;
   reg _392514_392514 ; 
   reg __392514_392514;
   reg _392515_392515 ; 
   reg __392515_392515;
   reg _392516_392516 ; 
   reg __392516_392516;
   reg _392517_392517 ; 
   reg __392517_392517;
   reg _392518_392518 ; 
   reg __392518_392518;
   reg _392519_392519 ; 
   reg __392519_392519;
   reg _392520_392520 ; 
   reg __392520_392520;
   reg _392521_392521 ; 
   reg __392521_392521;
   reg _392522_392522 ; 
   reg __392522_392522;
   reg _392523_392523 ; 
   reg __392523_392523;
   reg _392524_392524 ; 
   reg __392524_392524;
   reg _392525_392525 ; 
   reg __392525_392525;
   reg _392526_392526 ; 
   reg __392526_392526;
   reg _392527_392527 ; 
   reg __392527_392527;
   reg _392528_392528 ; 
   reg __392528_392528;
   reg _392529_392529 ; 
   reg __392529_392529;
   reg _392530_392530 ; 
   reg __392530_392530;
   reg _392531_392531 ; 
   reg __392531_392531;
   reg _392532_392532 ; 
   reg __392532_392532;
   reg _392533_392533 ; 
   reg __392533_392533;
   reg _392534_392534 ; 
   reg __392534_392534;
   reg _392535_392535 ; 
   reg __392535_392535;
   reg _392536_392536 ; 
   reg __392536_392536;
   reg _392537_392537 ; 
   reg __392537_392537;
   reg _392538_392538 ; 
   reg __392538_392538;
   reg _392539_392539 ; 
   reg __392539_392539;
   reg _392540_392540 ; 
   reg __392540_392540;
   reg _392541_392541 ; 
   reg __392541_392541;
   reg _392542_392542 ; 
   reg __392542_392542;
   reg _392543_392543 ; 
   reg __392543_392543;
   reg _392544_392544 ; 
   reg __392544_392544;
   reg _392545_392545 ; 
   reg __392545_392545;
   reg _392546_392546 ; 
   reg __392546_392546;
   reg _392547_392547 ; 
   reg __392547_392547;
   reg _392548_392548 ; 
   reg __392548_392548;
   reg _392549_392549 ; 
   reg __392549_392549;
   reg _392550_392550 ; 
   reg __392550_392550;
   reg _392551_392551 ; 
   reg __392551_392551;
   reg _392552_392552 ; 
   reg __392552_392552;
   reg _392553_392553 ; 
   reg __392553_392553;
   reg _392554_392554 ; 
   reg __392554_392554;
   reg _392555_392555 ; 
   reg __392555_392555;
   reg _392556_392556 ; 
   reg __392556_392556;
   reg _392557_392557 ; 
   reg __392557_392557;
   reg _392558_392558 ; 
   reg __392558_392558;
   reg _392559_392559 ; 
   reg __392559_392559;
   reg _392560_392560 ; 
   reg __392560_392560;
   reg _392561_392561 ; 
   reg __392561_392561;
   reg _392562_392562 ; 
   reg __392562_392562;
   reg _392563_392563 ; 
   reg __392563_392563;
   reg _392564_392564 ; 
   reg __392564_392564;
   reg _392565_392565 ; 
   reg __392565_392565;
   reg _392566_392566 ; 
   reg __392566_392566;
   reg _392567_392567 ; 
   reg __392567_392567;
   reg _392568_392568 ; 
   reg __392568_392568;
   reg _392569_392569 ; 
   reg __392569_392569;
   reg _392570_392570 ; 
   reg __392570_392570;
   reg _392571_392571 ; 
   reg __392571_392571;
   reg _392572_392572 ; 
   reg __392572_392572;
   reg _392573_392573 ; 
   reg __392573_392573;
   reg _392574_392574 ; 
   reg __392574_392574;
   reg _392575_392575 ; 
   reg __392575_392575;
   reg _392576_392576 ; 
   reg __392576_392576;
   reg _392577_392577 ; 
   reg __392577_392577;
   reg _392578_392578 ; 
   reg __392578_392578;
   reg _392579_392579 ; 
   reg __392579_392579;
   reg _392580_392580 ; 
   reg __392580_392580;
   reg _392581_392581 ; 
   reg __392581_392581;
   reg _392582_392582 ; 
   reg __392582_392582;
   reg _392583_392583 ; 
   reg __392583_392583;
   reg _392584_392584 ; 
   reg __392584_392584;
   reg _392585_392585 ; 
   reg __392585_392585;
   reg _392586_392586 ; 
   reg __392586_392586;
   reg _392587_392587 ; 
   reg __392587_392587;
   reg _392588_392588 ; 
   reg __392588_392588;
   reg _392589_392589 ; 
   reg __392589_392589;
   reg _392590_392590 ; 
   reg __392590_392590;
   reg _392591_392591 ; 
   reg __392591_392591;
   reg _392592_392592 ; 
   reg __392592_392592;
   reg _392593_392593 ; 
   reg __392593_392593;
   reg _392594_392594 ; 
   reg __392594_392594;
   reg _392595_392595 ; 
   reg __392595_392595;
   reg _392596_392596 ; 
   reg __392596_392596;
   reg _392597_392597 ; 
   reg __392597_392597;
   reg _392598_392598 ; 
   reg __392598_392598;
   reg _392599_392599 ; 
   reg __392599_392599;
   reg _392600_392600 ; 
   reg __392600_392600;
   reg _392601_392601 ; 
   reg __392601_392601;
   reg _392602_392602 ; 
   reg __392602_392602;
   reg _392603_392603 ; 
   reg __392603_392603;
   reg _392604_392604 ; 
   reg __392604_392604;
   reg _392605_392605 ; 
   reg __392605_392605;
   reg _392606_392606 ; 
   reg __392606_392606;
   reg _392607_392607 ; 
   reg __392607_392607;
   reg _392608_392608 ; 
   reg __392608_392608;
   reg _392609_392609 ; 
   reg __392609_392609;
   reg _392610_392610 ; 
   reg __392610_392610;
   reg _392611_392611 ; 
   reg __392611_392611;
   reg _392612_392612 ; 
   reg __392612_392612;
   reg _392613_392613 ; 
   reg __392613_392613;
   reg _392614_392614 ; 
   reg __392614_392614;
   reg _392615_392615 ; 
   reg __392615_392615;
   reg _392616_392616 ; 
   reg __392616_392616;
   reg _392617_392617 ; 
   reg __392617_392617;
   reg _392618_392618 ; 
   reg __392618_392618;
   reg _392619_392619 ; 
   reg __392619_392619;
   reg _392620_392620 ; 
   reg __392620_392620;
   reg _392621_392621 ; 
   reg __392621_392621;
   reg _392622_392622 ; 
   reg __392622_392622;
   reg _392623_392623 ; 
   reg __392623_392623;
   reg _392624_392624 ; 
   reg __392624_392624;
   reg _392625_392625 ; 
   reg __392625_392625;
   reg _392626_392626 ; 
   reg __392626_392626;
   reg _392627_392627 ; 
   reg __392627_392627;
   reg _392628_392628 ; 
   reg __392628_392628;
   reg _392629_392629 ; 
   reg __392629_392629;
   reg _392630_392630 ; 
   reg __392630_392630;
   reg _392631_392631 ; 
   reg __392631_392631;
   reg _392632_392632 ; 
   reg __392632_392632;
   reg _392633_392633 ; 
   reg __392633_392633;
   reg _392634_392634 ; 
   reg __392634_392634;
   reg _392635_392635 ; 
   reg __392635_392635;
   reg _392636_392636 ; 
   reg __392636_392636;
   reg _392637_392637 ; 
   reg __392637_392637;
   reg _392638_392638 ; 
   reg __392638_392638;
   reg _392639_392639 ; 
   reg __392639_392639;
   reg _392640_392640 ; 
   reg __392640_392640;
   reg _392641_392641 ; 
   reg __392641_392641;
   reg _392642_392642 ; 
   reg __392642_392642;
   reg _392643_392643 ; 
   reg __392643_392643;
   reg _392644_392644 ; 
   reg __392644_392644;
   reg _392645_392645 ; 
   reg __392645_392645;
   reg _392646_392646 ; 
   reg __392646_392646;
   reg _392647_392647 ; 
   reg __392647_392647;
   reg _392648_392648 ; 
   reg __392648_392648;
   reg _392649_392649 ; 
   reg __392649_392649;
   reg _392650_392650 ; 
   reg __392650_392650;
   reg _392651_392651 ; 
   reg __392651_392651;
   reg _392652_392652 ; 
   reg __392652_392652;
   reg _392653_392653 ; 
   reg __392653_392653;
   reg _392654_392654 ; 
   reg __392654_392654;
   reg _392655_392655 ; 
   reg __392655_392655;
   reg _392656_392656 ; 
   reg __392656_392656;
   reg _392657_392657 ; 
   reg __392657_392657;
   reg _392658_392658 ; 
   reg __392658_392658;
   reg _392659_392659 ; 
   reg __392659_392659;
   reg _392660_392660 ; 
   reg __392660_392660;
   reg _392661_392661 ; 
   reg __392661_392661;
   reg _392662_392662 ; 
   reg __392662_392662;
   reg _392663_392663 ; 
   reg __392663_392663;
   reg _392664_392664 ; 
   reg __392664_392664;
   reg _392665_392665 ; 
   reg __392665_392665;
   reg _392666_392666 ; 
   reg __392666_392666;
   reg _392667_392667 ; 
   reg __392667_392667;
   reg _392668_392668 ; 
   reg __392668_392668;
   reg _392669_392669 ; 
   reg __392669_392669;
   reg _392670_392670 ; 
   reg __392670_392670;
   reg _392671_392671 ; 
   reg __392671_392671;
   reg _392672_392672 ; 
   reg __392672_392672;
   reg _392673_392673 ; 
   reg __392673_392673;
   reg _392674_392674 ; 
   reg __392674_392674;
   reg _392675_392675 ; 
   reg __392675_392675;
   reg _392676_392676 ; 
   reg __392676_392676;
   reg _392677_392677 ; 
   reg __392677_392677;
   reg _392678_392678 ; 
   reg __392678_392678;
   reg _392679_392679 ; 
   reg __392679_392679;
   reg _392680_392680 ; 
   reg __392680_392680;
   reg _392681_392681 ; 
   reg __392681_392681;
   reg _392682_392682 ; 
   reg __392682_392682;
   reg _392683_392683 ; 
   reg __392683_392683;
   reg _392684_392684 ; 
   reg __392684_392684;
   reg _392685_392685 ; 
   reg __392685_392685;
   reg _392686_392686 ; 
   reg __392686_392686;
   reg _392687_392687 ; 
   reg __392687_392687;
   reg _392688_392688 ; 
   reg __392688_392688;
   reg _392689_392689 ; 
   reg __392689_392689;
   reg _392690_392690 ; 
   reg __392690_392690;
   reg _392691_392691 ; 
   reg __392691_392691;
   reg _392692_392692 ; 
   reg __392692_392692;
   reg _392693_392693 ; 
   reg __392693_392693;
   reg _392694_392694 ; 
   reg __392694_392694;
   reg _392695_392695 ; 
   reg __392695_392695;
   reg _392696_392696 ; 
   reg __392696_392696;
   reg _392697_392697 ; 
   reg __392697_392697;
   reg _392698_392698 ; 
   reg __392698_392698;
   reg _392699_392699 ; 
   reg __392699_392699;
   reg _392700_392700 ; 
   reg __392700_392700;
   reg _392701_392701 ; 
   reg __392701_392701;
   reg _392702_392702 ; 
   reg __392702_392702;
   reg _392703_392703 ; 
   reg __392703_392703;
   reg _392704_392704 ; 
   reg __392704_392704;
   reg _392705_392705 ; 
   reg __392705_392705;
   reg _392706_392706 ; 
   reg __392706_392706;
   reg _392707_392707 ; 
   reg __392707_392707;
   reg _392708_392708 ; 
   reg __392708_392708;
   reg _392709_392709 ; 
   reg __392709_392709;
   reg _392710_392710 ; 
   reg __392710_392710;
   reg _392711_392711 ; 
   reg __392711_392711;
   reg _392712_392712 ; 
   reg __392712_392712;
   reg _392713_392713 ; 
   reg __392713_392713;
   reg _392714_392714 ; 
   reg __392714_392714;
   reg _392715_392715 ; 
   reg __392715_392715;
   reg _392716_392716 ; 
   reg __392716_392716;
   reg _392717_392717 ; 
   reg __392717_392717;
   reg _392718_392718 ; 
   reg __392718_392718;
   reg _392719_392719 ; 
   reg __392719_392719;
   reg _392720_392720 ; 
   reg __392720_392720;
   reg _392721_392721 ; 
   reg __392721_392721;
   reg _392722_392722 ; 
   reg __392722_392722;
   reg _392723_392723 ; 
   reg __392723_392723;
   reg _392724_392724 ; 
   reg __392724_392724;
   reg _392725_392725 ; 
   reg __392725_392725;
   reg _392726_392726 ; 
   reg __392726_392726;
   reg _392727_392727 ; 
   reg __392727_392727;
   reg _392728_392728 ; 
   reg __392728_392728;
   reg _392729_392729 ; 
   reg __392729_392729;
   reg _392730_392730 ; 
   reg __392730_392730;
   reg _392731_392731 ; 
   reg __392731_392731;
   reg _392732_392732 ; 
   reg __392732_392732;
   reg _392733_392733 ; 
   reg __392733_392733;
   reg _392734_392734 ; 
   reg __392734_392734;
   reg _392735_392735 ; 
   reg __392735_392735;
   reg _392736_392736 ; 
   reg __392736_392736;
   reg _392737_392737 ; 
   reg __392737_392737;
   reg _392738_392738 ; 
   reg __392738_392738;
   reg _392739_392739 ; 
   reg __392739_392739;
   reg _392740_392740 ; 
   reg __392740_392740;
   reg _392741_392741 ; 
   reg __392741_392741;
   reg _392742_392742 ; 
   reg __392742_392742;
   reg _392743_392743 ; 
   reg __392743_392743;
   reg _392744_392744 ; 
   reg __392744_392744;
   reg _392745_392745 ; 
   reg __392745_392745;
   reg _392746_392746 ; 
   reg __392746_392746;
   reg _392747_392747 ; 
   reg __392747_392747;
   reg _392748_392748 ; 
   reg __392748_392748;
   reg _392749_392749 ; 
   reg __392749_392749;
   reg _392750_392750 ; 
   reg __392750_392750;
   reg _392751_392751 ; 
   reg __392751_392751;
   reg _392752_392752 ; 
   reg __392752_392752;
   reg _392753_392753 ; 
   reg __392753_392753;
   reg _392754_392754 ; 
   reg __392754_392754;
   reg _392755_392755 ; 
   reg __392755_392755;
   reg _392756_392756 ; 
   reg __392756_392756;
   reg _392757_392757 ; 
   reg __392757_392757;
   reg _392758_392758 ; 
   reg __392758_392758;
   reg _392759_392759 ; 
   reg __392759_392759;
   reg _392760_392760 ; 
   reg __392760_392760;
   reg _392761_392761 ; 
   reg __392761_392761;
   reg _392762_392762 ; 
   reg __392762_392762;
   reg _392763_392763 ; 
   reg __392763_392763;
   reg _392764_392764 ; 
   reg __392764_392764;
   reg _392765_392765 ; 
   reg __392765_392765;
   reg _392766_392766 ; 
   reg __392766_392766;
   reg _392767_392767 ; 
   reg __392767_392767;
   reg _392768_392768 ; 
   reg __392768_392768;
   reg _392769_392769 ; 
   reg __392769_392769;
   reg _392770_392770 ; 
   reg __392770_392770;
   reg _392771_392771 ; 
   reg __392771_392771;
   reg _392772_392772 ; 
   reg __392772_392772;
   reg _392773_392773 ; 
   reg __392773_392773;
   reg _392774_392774 ; 
   reg __392774_392774;
   reg _392775_392775 ; 
   reg __392775_392775;
   reg _392776_392776 ; 
   reg __392776_392776;
   reg _392777_392777 ; 
   reg __392777_392777;
   reg _392778_392778 ; 
   reg __392778_392778;
   reg _392779_392779 ; 
   reg __392779_392779;
   reg _392780_392780 ; 
   reg __392780_392780;
   reg _392781_392781 ; 
   reg __392781_392781;
   reg _392782_392782 ; 
   reg __392782_392782;
   reg _392783_392783 ; 
   reg __392783_392783;
   reg _392784_392784 ; 
   reg __392784_392784;
   reg _392785_392785 ; 
   reg __392785_392785;
   reg _392786_392786 ; 
   reg __392786_392786;
   reg _392787_392787 ; 
   reg __392787_392787;
   reg _392788_392788 ; 
   reg __392788_392788;
   reg _392789_392789 ; 
   reg __392789_392789;
   reg _392790_392790 ; 
   reg __392790_392790;
   reg _392791_392791 ; 
   reg __392791_392791;
   reg _392792_392792 ; 
   reg __392792_392792;
   reg _392793_392793 ; 
   reg __392793_392793;
   reg _392794_392794 ; 
   reg __392794_392794;
   reg _392795_392795 ; 
   reg __392795_392795;
   reg _392796_392796 ; 
   reg __392796_392796;
   reg _392797_392797 ; 
   reg __392797_392797;
   reg _392798_392798 ; 
   reg __392798_392798;
   reg _392799_392799 ; 
   reg __392799_392799;
   reg _392800_392800 ; 
   reg __392800_392800;
   reg _392801_392801 ; 
   reg __392801_392801;
   reg _392802_392802 ; 
   reg __392802_392802;
   reg _392803_392803 ; 
   reg __392803_392803;
   reg _392804_392804 ; 
   reg __392804_392804;
   reg _392805_392805 ; 
   reg __392805_392805;
   reg _392806_392806 ; 
   reg __392806_392806;
   reg _392807_392807 ; 
   reg __392807_392807;
   reg _392808_392808 ; 
   reg __392808_392808;
   reg _392809_392809 ; 
   reg __392809_392809;
   reg _392810_392810 ; 
   reg __392810_392810;
   reg _392811_392811 ; 
   reg __392811_392811;
   reg _392812_392812 ; 
   reg __392812_392812;
   reg _392813_392813 ; 
   reg __392813_392813;
   reg _392814_392814 ; 
   reg __392814_392814;
   reg _392815_392815 ; 
   reg __392815_392815;
   reg _392816_392816 ; 
   reg __392816_392816;
   reg _392817_392817 ; 
   reg __392817_392817;
   reg _392818_392818 ; 
   reg __392818_392818;
   reg _392819_392819 ; 
   reg __392819_392819;
   reg _392820_392820 ; 
   reg __392820_392820;
   reg _392821_392821 ; 
   reg __392821_392821;
   reg _392822_392822 ; 
   reg __392822_392822;
   reg _392823_392823 ; 
   reg __392823_392823;
   reg _392824_392824 ; 
   reg __392824_392824;
   reg _392825_392825 ; 
   reg __392825_392825;
   reg _392826_392826 ; 
   reg __392826_392826;
   reg _392827_392827 ; 
   reg __392827_392827;
   reg _392828_392828 ; 
   reg __392828_392828;
   reg _392829_392829 ; 
   reg __392829_392829;
   reg _392830_392830 ; 
   reg __392830_392830;
   reg _392831_392831 ; 
   reg __392831_392831;
   reg _392832_392832 ; 
   reg __392832_392832;
   reg _392833_392833 ; 
   reg __392833_392833;
   reg _392834_392834 ; 
   reg __392834_392834;
   reg _392835_392835 ; 
   reg __392835_392835;
   reg _392836_392836 ; 
   reg __392836_392836;
   reg _392837_392837 ; 
   reg __392837_392837;
   reg _392838_392838 ; 
   reg __392838_392838;
   reg _392839_392839 ; 
   reg __392839_392839;
   reg _392840_392840 ; 
   reg __392840_392840;
   reg _392841_392841 ; 
   reg __392841_392841;
   reg _392842_392842 ; 
   reg __392842_392842;
   reg _392843_392843 ; 
   reg __392843_392843;
   reg _392844_392844 ; 
   reg __392844_392844;
   reg _392845_392845 ; 
   reg __392845_392845;
   reg _392846_392846 ; 
   reg __392846_392846;
   reg _392847_392847 ; 
   reg __392847_392847;
   reg _392848_392848 ; 
   reg __392848_392848;
   reg _392849_392849 ; 
   reg __392849_392849;
   reg _392850_392850 ; 
   reg __392850_392850;
   reg _392851_392851 ; 
   reg __392851_392851;
   reg _392852_392852 ; 
   reg __392852_392852;
   reg _392853_392853 ; 
   reg __392853_392853;
   reg _392854_392854 ; 
   reg __392854_392854;
   reg _392855_392855 ; 
   reg __392855_392855;
   reg _392856_392856 ; 
   reg __392856_392856;
   reg _392857_392857 ; 
   reg __392857_392857;
   reg _392858_392858 ; 
   reg __392858_392858;
   reg _392859_392859 ; 
   reg __392859_392859;
   reg _392860_392860 ; 
   reg __392860_392860;
   reg _392861_392861 ; 
   reg __392861_392861;
   reg _392862_392862 ; 
   reg __392862_392862;
   reg _392863_392863 ; 
   reg __392863_392863;
   reg _392864_392864 ; 
   reg __392864_392864;
   reg _392865_392865 ; 
   reg __392865_392865;
   reg _392866_392866 ; 
   reg __392866_392866;
   reg _392867_392867 ; 
   reg __392867_392867;
   reg _392868_392868 ; 
   reg __392868_392868;
   reg _392869_392869 ; 
   reg __392869_392869;
   reg _392870_392870 ; 
   reg __392870_392870;
   reg _392871_392871 ; 
   reg __392871_392871;
   reg _392872_392872 ; 
   reg __392872_392872;
   reg _392873_392873 ; 
   reg __392873_392873;
   reg _392874_392874 ; 
   reg __392874_392874;
   reg _392875_392875 ; 
   reg __392875_392875;
   reg _392876_392876 ; 
   reg __392876_392876;
   reg _392877_392877 ; 
   reg __392877_392877;
   reg _392878_392878 ; 
   reg __392878_392878;
   reg _392879_392879 ; 
   reg __392879_392879;
   reg _392880_392880 ; 
   reg __392880_392880;
   reg _392881_392881 ; 
   reg __392881_392881;
   reg _392882_392882 ; 
   reg __392882_392882;
   reg _392883_392883 ; 
   reg __392883_392883;
   reg _392884_392884 ; 
   reg __392884_392884;
   reg _392885_392885 ; 
   reg __392885_392885;
   reg _392886_392886 ; 
   reg __392886_392886;
   reg _392887_392887 ; 
   reg __392887_392887;
   reg _392888_392888 ; 
   reg __392888_392888;
   reg _392889_392889 ; 
   reg __392889_392889;
   reg _392890_392890 ; 
   reg __392890_392890;
   reg _392891_392891 ; 
   reg __392891_392891;
   reg _392892_392892 ; 
   reg __392892_392892;
   reg _392893_392893 ; 
   reg __392893_392893;
   reg _392894_392894 ; 
   reg __392894_392894;
   reg _392895_392895 ; 
   reg __392895_392895;
   reg _392896_392896 ; 
   reg __392896_392896;
   reg _392897_392897 ; 
   reg __392897_392897;
   reg _392898_392898 ; 
   reg __392898_392898;
   reg _392899_392899 ; 
   reg __392899_392899;
   reg _392900_392900 ; 
   reg __392900_392900;
   reg _392901_392901 ; 
   reg __392901_392901;
   reg _392902_392902 ; 
   reg __392902_392902;
   reg _392903_392903 ; 
   reg __392903_392903;
   reg _392904_392904 ; 
   reg __392904_392904;
   reg _392905_392905 ; 
   reg __392905_392905;
   reg _392906_392906 ; 
   reg __392906_392906;
   reg _392907_392907 ; 
   reg __392907_392907;
   reg _392908_392908 ; 
   reg __392908_392908;
   reg _392909_392909 ; 
   reg __392909_392909;
   reg _392910_392910 ; 
   reg __392910_392910;
   reg _392911_392911 ; 
   reg __392911_392911;
   reg _392912_392912 ; 
   reg __392912_392912;
   reg _392913_392913 ; 
   reg __392913_392913;
   reg _392914_392914 ; 
   reg __392914_392914;
   reg _392915_392915 ; 
   reg __392915_392915;
   reg _392916_392916 ; 
   reg __392916_392916;
   reg _392917_392917 ; 
   reg __392917_392917;
   reg _392918_392918 ; 
   reg __392918_392918;
   reg _392919_392919 ; 
   reg __392919_392919;
   reg _392920_392920 ; 
   reg __392920_392920;
   reg _392921_392921 ; 
   reg __392921_392921;
   reg _392922_392922 ; 
   reg __392922_392922;
   reg _392923_392923 ; 
   reg __392923_392923;
   reg _392924_392924 ; 
   reg __392924_392924;
   reg _392925_392925 ; 
   reg __392925_392925;
   reg _392926_392926 ; 
   reg __392926_392926;
   reg _392927_392927 ; 
   reg __392927_392927;
   reg _392928_392928 ; 
   reg __392928_392928;
   reg _392929_392929 ; 
   reg __392929_392929;
   reg _392930_392930 ; 
   reg __392930_392930;
   reg _392931_392931 ; 
   reg __392931_392931;
   reg _392932_392932 ; 
   reg __392932_392932;
   reg _392933_392933 ; 
   reg __392933_392933;
   reg _392934_392934 ; 
   reg __392934_392934;
   reg _392935_392935 ; 
   reg __392935_392935;
   reg _392936_392936 ; 
   reg __392936_392936;
   reg _392937_392937 ; 
   reg __392937_392937;
   reg _392938_392938 ; 
   reg __392938_392938;
   reg _392939_392939 ; 
   reg __392939_392939;
   reg _392940_392940 ; 
   reg __392940_392940;
   reg _392941_392941 ; 
   reg __392941_392941;
   reg _392942_392942 ; 
   reg __392942_392942;
   reg _392943_392943 ; 
   reg __392943_392943;
   reg _392944_392944 ; 
   reg __392944_392944;
   reg _392945_392945 ; 
   reg __392945_392945;
   reg _392946_392946 ; 
   reg __392946_392946;
   reg _392947_392947 ; 
   reg __392947_392947;
   reg _392948_392948 ; 
   reg __392948_392948;
   reg _392949_392949 ; 
   reg __392949_392949;
   reg _392950_392950 ; 
   reg __392950_392950;
   reg _392951_392951 ; 
   reg __392951_392951;
   reg _392952_392952 ; 
   reg __392952_392952;
   reg _392953_392953 ; 
   reg __392953_392953;
   reg _392954_392954 ; 
   reg __392954_392954;
   reg _392955_392955 ; 
   reg __392955_392955;
   reg _392956_392956 ; 
   reg __392956_392956;
   reg _392957_392957 ; 
   reg __392957_392957;
   reg _392958_392958 ; 
   reg __392958_392958;
   reg _392959_392959 ; 
   reg __392959_392959;
   reg _392960_392960 ; 
   reg __392960_392960;
   reg _392961_392961 ; 
   reg __392961_392961;
   reg _392962_392962 ; 
   reg __392962_392962;
   reg _392963_392963 ; 
   reg __392963_392963;
   reg _392964_392964 ; 
   reg __392964_392964;
   reg _392965_392965 ; 
   reg __392965_392965;
   reg _392966_392966 ; 
   reg __392966_392966;
   reg _392967_392967 ; 
   reg __392967_392967;
   reg _392968_392968 ; 
   reg __392968_392968;
   reg _392969_392969 ; 
   reg __392969_392969;
   reg _392970_392970 ; 
   reg __392970_392970;
   reg _392971_392971 ; 
   reg __392971_392971;
   reg _392972_392972 ; 
   reg __392972_392972;
   reg _392973_392973 ; 
   reg __392973_392973;
   reg _392974_392974 ; 
   reg __392974_392974;
   reg _392975_392975 ; 
   reg __392975_392975;
   reg _392976_392976 ; 
   reg __392976_392976;
   reg _392977_392977 ; 
   reg __392977_392977;
   reg _392978_392978 ; 
   reg __392978_392978;
   reg _392979_392979 ; 
   reg __392979_392979;
   reg _392980_392980 ; 
   reg __392980_392980;
   reg _392981_392981 ; 
   reg __392981_392981;
   reg _392982_392982 ; 
   reg __392982_392982;
   reg _392983_392983 ; 
   reg __392983_392983;
   reg _392984_392984 ; 
   reg __392984_392984;
   reg _392985_392985 ; 
   reg __392985_392985;
   reg _392986_392986 ; 
   reg __392986_392986;
   reg _392987_392987 ; 
   reg __392987_392987;
   reg _392988_392988 ; 
   reg __392988_392988;
   reg _392989_392989 ; 
   reg __392989_392989;
   reg _392990_392990 ; 
   reg __392990_392990;
   reg _392991_392991 ; 
   reg __392991_392991;
   reg _392992_392992 ; 
   reg __392992_392992;
   reg _392993_392993 ; 
   reg __392993_392993;
   reg _392994_392994 ; 
   reg __392994_392994;
   reg _392995_392995 ; 
   reg __392995_392995;
   reg _392996_392996 ; 
   reg __392996_392996;
   reg _392997_392997 ; 
   reg __392997_392997;
   reg _392998_392998 ; 
   reg __392998_392998;
   reg _392999_392999 ; 
   reg __392999_392999;
   reg _393000_393000 ; 
   reg __393000_393000;
   reg _393001_393001 ; 
   reg __393001_393001;
   reg _393002_393002 ; 
   reg __393002_393002;
   reg _393003_393003 ; 
   reg __393003_393003;
   reg _393004_393004 ; 
   reg __393004_393004;
   reg _393005_393005 ; 
   reg __393005_393005;
   reg _393006_393006 ; 
   reg __393006_393006;
   reg _393007_393007 ; 
   reg __393007_393007;
   reg _393008_393008 ; 
   reg __393008_393008;
   reg _393009_393009 ; 
   reg __393009_393009;
   reg _393010_393010 ; 
   reg __393010_393010;
   reg _393011_393011 ; 
   reg __393011_393011;
   reg _393012_393012 ; 
   reg __393012_393012;
   reg _393013_393013 ; 
   reg __393013_393013;
   reg _393014_393014 ; 
   reg __393014_393014;
   reg _393015_393015 ; 
   reg __393015_393015;
   reg _393016_393016 ; 
   reg __393016_393016;
   reg _393017_393017 ; 
   reg __393017_393017;
   reg _393018_393018 ; 
   reg __393018_393018;
   reg _393019_393019 ; 
   reg __393019_393019;
   reg _393020_393020 ; 
   reg __393020_393020;
   reg _393021_393021 ; 
   reg __393021_393021;
   reg _393022_393022 ; 
   reg __393022_393022;
   reg _393023_393023 ; 
   reg __393023_393023;
   reg _393024_393024 ; 
   reg __393024_393024;
   reg _393025_393025 ; 
   reg __393025_393025;
   reg _393026_393026 ; 
   reg __393026_393026;
   reg _393027_393027 ; 
   reg __393027_393027;
   reg _393028_393028 ; 
   reg __393028_393028;
   reg _393029_393029 ; 
   reg __393029_393029;
   reg _393030_393030 ; 
   reg __393030_393030;
   reg _393031_393031 ; 
   reg __393031_393031;
   reg _393032_393032 ; 
   reg __393032_393032;
   reg _393033_393033 ; 
   reg __393033_393033;
   reg _393034_393034 ; 
   reg __393034_393034;
   reg _393035_393035 ; 
   reg __393035_393035;
   reg _393036_393036 ; 
   reg __393036_393036;
   reg _393037_393037 ; 
   reg __393037_393037;
   reg _393038_393038 ; 
   reg __393038_393038;
   reg _393039_393039 ; 
   reg __393039_393039;
   reg _393040_393040 ; 
   reg __393040_393040;
   reg _393041_393041 ; 
   reg __393041_393041;
   reg _393042_393042 ; 
   reg __393042_393042;
   reg _393043_393043 ; 
   reg __393043_393043;
   reg _393044_393044 ; 
   reg __393044_393044;
   reg _393045_393045 ; 
   reg __393045_393045;
   reg _393046_393046 ; 
   reg __393046_393046;
   reg _393047_393047 ; 
   reg __393047_393047;
   reg _393048_393048 ; 
   reg __393048_393048;
   reg _393049_393049 ; 
   reg __393049_393049;
   reg _393050_393050 ; 
   reg __393050_393050;
   reg _393051_393051 ; 
   reg __393051_393051;
   reg _393052_393052 ; 
   reg __393052_393052;
   reg _393053_393053 ; 
   reg __393053_393053;
   reg _393054_393054 ; 
   reg __393054_393054;
   reg _393055_393055 ; 
   reg __393055_393055;
   reg _393056_393056 ; 
   reg __393056_393056;
   reg _393057_393057 ; 
   reg __393057_393057;
   reg _393058_393058 ; 
   reg __393058_393058;
   reg _393059_393059 ; 
   reg __393059_393059;
   reg _393060_393060 ; 
   reg __393060_393060;
   reg _393061_393061 ; 
   reg __393061_393061;
   reg _393062_393062 ; 
   reg __393062_393062;
   reg _393063_393063 ; 
   reg __393063_393063;
   reg _393064_393064 ; 
   reg __393064_393064;
   reg _393065_393065 ; 
   reg __393065_393065;
   reg _393066_393066 ; 
   reg __393066_393066;
   reg _393067_393067 ; 
   reg __393067_393067;
   reg _393068_393068 ; 
   reg __393068_393068;
   reg _393069_393069 ; 
   reg __393069_393069;
   reg _393070_393070 ; 
   reg __393070_393070;
   reg _393071_393071 ; 
   reg __393071_393071;
   reg _393072_393072 ; 
   reg __393072_393072;
   reg _393073_393073 ; 
   reg __393073_393073;
   reg _393074_393074 ; 
   reg __393074_393074;
   reg _393075_393075 ; 
   reg __393075_393075;
   reg _393076_393076 ; 
   reg __393076_393076;
   reg _393077_393077 ; 
   reg __393077_393077;
   reg _393078_393078 ; 
   reg __393078_393078;
   reg _393079_393079 ; 
   reg __393079_393079;
   reg _393080_393080 ; 
   reg __393080_393080;
   reg _393081_393081 ; 
   reg __393081_393081;
   reg _393082_393082 ; 
   reg __393082_393082;
   reg _393083_393083 ; 
   reg __393083_393083;
   reg _393084_393084 ; 
   reg __393084_393084;
   reg _393085_393085 ; 
   reg __393085_393085;
   reg _393086_393086 ; 
   reg __393086_393086;
   reg _393087_393087 ; 
   reg __393087_393087;
   reg _393088_393088 ; 
   reg __393088_393088;
   reg _393089_393089 ; 
   reg __393089_393089;
   reg _393090_393090 ; 
   reg __393090_393090;
   reg _393091_393091 ; 
   reg __393091_393091;
   reg _393092_393092 ; 
   reg __393092_393092;
   reg _393093_393093 ; 
   reg __393093_393093;
   reg _393094_393094 ; 
   reg __393094_393094;
   reg _393095_393095 ; 
   reg __393095_393095;
   reg _393096_393096 ; 
   reg __393096_393096;
   reg _393097_393097 ; 
   reg __393097_393097;
   reg _393098_393098 ; 
   reg __393098_393098;
   reg _393099_393099 ; 
   reg __393099_393099;
   reg _393100_393100 ; 
   reg __393100_393100;
   reg _393101_393101 ; 
   reg __393101_393101;
   reg _393102_393102 ; 
   reg __393102_393102;
   reg _393103_393103 ; 
   reg __393103_393103;
   reg _393104_393104 ; 
   reg __393104_393104;
   reg _393105_393105 ; 
   reg __393105_393105;
   reg _393106_393106 ; 
   reg __393106_393106;
   reg _393107_393107 ; 
   reg __393107_393107;
   reg _393108_393108 ; 
   reg __393108_393108;
   reg _393109_393109 ; 
   reg __393109_393109;
   reg _393110_393110 ; 
   reg __393110_393110;
   reg _393111_393111 ; 
   reg __393111_393111;
   reg _393112_393112 ; 
   reg __393112_393112;
   reg _393113_393113 ; 
   reg __393113_393113;
   reg _393114_393114 ; 
   reg __393114_393114;
   reg _393115_393115 ; 
   reg __393115_393115;
   reg _393116_393116 ; 
   reg __393116_393116;
   reg _393117_393117 ; 
   reg __393117_393117;
   reg _393118_393118 ; 
   reg __393118_393118;
   reg _393119_393119 ; 
   reg __393119_393119;
   reg _393120_393120 ; 
   reg __393120_393120;
   reg _393121_393121 ; 
   reg __393121_393121;
   reg _393122_393122 ; 
   reg __393122_393122;
   reg _393123_393123 ; 
   reg __393123_393123;
   reg _393124_393124 ; 
   reg __393124_393124;
   reg _393125_393125 ; 
   reg __393125_393125;
   reg _393126_393126 ; 
   reg __393126_393126;
   reg _393127_393127 ; 
   reg __393127_393127;
   reg _393128_393128 ; 
   reg __393128_393128;
   reg _393129_393129 ; 
   reg __393129_393129;
   reg _393130_393130 ; 
   reg __393130_393130;
   reg _393131_393131 ; 
   reg __393131_393131;
   reg _393132_393132 ; 
   reg __393132_393132;
   reg _393133_393133 ; 
   reg __393133_393133;
   reg _393134_393134 ; 
   reg __393134_393134;
   reg _393135_393135 ; 
   reg __393135_393135;
   reg _393136_393136 ; 
   reg __393136_393136;
   reg _393137_393137 ; 
   reg __393137_393137;
   reg _393138_393138 ; 
   reg __393138_393138;
   reg _393139_393139 ; 
   reg __393139_393139;
   reg _393140_393140 ; 
   reg __393140_393140;
   reg _393141_393141 ; 
   reg __393141_393141;
   reg _393142_393142 ; 
   reg __393142_393142;
   reg _393143_393143 ; 
   reg __393143_393143;
   reg _393144_393144 ; 
   reg __393144_393144;
   reg _393145_393145 ; 
   reg __393145_393145;
   reg _393146_393146 ; 
   reg __393146_393146;
   reg _393147_393147 ; 
   reg __393147_393147;
   reg _393148_393148 ; 
   reg __393148_393148;
   reg _393149_393149 ; 
   reg __393149_393149;
   reg _393150_393150 ; 
   reg __393150_393150;
   reg _393151_393151 ; 
   reg __393151_393151;
   reg _393152_393152 ; 
   reg __393152_393152;
   reg _393153_393153 ; 
   reg __393153_393153;
   reg _393154_393154 ; 
   reg __393154_393154;
   reg _393155_393155 ; 
   reg __393155_393155;
   reg _393156_393156 ; 
   reg __393156_393156;
   reg _393157_393157 ; 
   reg __393157_393157;
   reg _393158_393158 ; 
   reg __393158_393158;
   reg _393159_393159 ; 
   reg __393159_393159;
   reg _393160_393160 ; 
   reg __393160_393160;
   reg _393161_393161 ; 
   reg __393161_393161;
   reg _393162_393162 ; 
   reg __393162_393162;
   reg _393163_393163 ; 
   reg __393163_393163;
   reg _393164_393164 ; 
   reg __393164_393164;
   reg _393165_393165 ; 
   reg __393165_393165;
   reg _393166_393166 ; 
   reg __393166_393166;
   reg _393167_393167 ; 
   reg __393167_393167;
   reg _393168_393168 ; 
   reg __393168_393168;
   reg _393169_393169 ; 
   reg __393169_393169;
   reg _393170_393170 ; 
   reg __393170_393170;
   reg _393171_393171 ; 
   reg __393171_393171;
   reg _393172_393172 ; 
   reg __393172_393172;
   reg _393173_393173 ; 
   reg __393173_393173;
   reg _393174_393174 ; 
   reg __393174_393174;
   reg _393175_393175 ; 
   reg __393175_393175;
   reg _393176_393176 ; 
   reg __393176_393176;
   reg _393177_393177 ; 
   reg __393177_393177;
   reg _393178_393178 ; 
   reg __393178_393178;
   reg _393179_393179 ; 
   reg __393179_393179;
   reg _393180_393180 ; 
   reg __393180_393180;
   reg _393181_393181 ; 
   reg __393181_393181;
   reg _393182_393182 ; 
   reg __393182_393182;
   reg _393183_393183 ; 
   reg __393183_393183;
   reg _393184_393184 ; 
   reg __393184_393184;
   reg _393185_393185 ; 
   reg __393185_393185;
   reg _393186_393186 ; 
   reg __393186_393186;
   reg _393187_393187 ; 
   reg __393187_393187;
   reg _393188_393188 ; 
   reg __393188_393188;
   reg _393189_393189 ; 
   reg __393189_393189;
   reg _393190_393190 ; 
   reg __393190_393190;
   reg _393191_393191 ; 
   reg __393191_393191;
   reg _393192_393192 ; 
   reg __393192_393192;
   reg _393193_393193 ; 
   reg __393193_393193;
   reg _393194_393194 ; 
   reg __393194_393194;
   reg _393195_393195 ; 
   reg __393195_393195;
   reg _393196_393196 ; 
   reg __393196_393196;
   reg _393197_393197 ; 
   reg __393197_393197;
   reg _393198_393198 ; 
   reg __393198_393198;
   reg _393199_393199 ; 
   reg __393199_393199;
   reg _393200_393200 ; 
   reg __393200_393200;
   reg _393201_393201 ; 
   reg __393201_393201;
   reg _393202_393202 ; 
   reg __393202_393202;
   reg _393203_393203 ; 
   reg __393203_393203;
   reg _393204_393204 ; 
   reg __393204_393204;
   reg _393205_393205 ; 
   reg __393205_393205;
   reg _393206_393206 ; 
   reg __393206_393206;
   reg _393207_393207 ; 
   reg __393207_393207;
   reg _393208_393208 ; 
   reg __393208_393208;
   reg _393209_393209 ; 
   reg __393209_393209;
   reg _393210_393210 ; 
   reg __393210_393210;
   reg _393211_393211 ; 
   reg __393211_393211;
   reg _393212_393212 ; 
   reg __393212_393212;
   reg _393213_393213 ; 
   reg __393213_393213;
   reg _393214_393214 ; 
   reg __393214_393214;
   reg _393215_393215 ; 
   reg __393215_393215;
   reg _393216_393216 ; 
   reg __393216_393216;
   reg _393217_393217 ; 
   reg __393217_393217;
   reg _393218_393218 ; 
   reg __393218_393218;
   reg _393219_393219 ; 
   reg __393219_393219;
   reg _393220_393220 ; 
   reg __393220_393220;
   reg _393221_393221 ; 
   reg __393221_393221;
   reg _393222_393222 ; 
   reg __393222_393222;
   reg _393223_393223 ; 
   reg __393223_393223;
   reg _393224_393224 ; 
   reg __393224_393224;
   reg _393225_393225 ; 
   reg __393225_393225;
   reg _393226_393226 ; 
   reg __393226_393226;
   reg _393227_393227 ; 
   reg __393227_393227;
   reg _393228_393228 ; 
   reg __393228_393228;
   reg _393229_393229 ; 
   reg __393229_393229;
   reg _393230_393230 ; 
   reg __393230_393230;
   reg _393231_393231 ; 
   reg __393231_393231;
   reg _393232_393232 ; 
   reg __393232_393232;
   reg _393233_393233 ; 
   reg __393233_393233;
   reg _393234_393234 ; 
   reg __393234_393234;
   reg _393235_393235 ; 
   reg __393235_393235;
   reg _393236_393236 ; 
   reg __393236_393236;
   reg _393237_393237 ; 
   reg __393237_393237;
   reg _393238_393238 ; 
   reg __393238_393238;
   reg _393239_393239 ; 
   reg __393239_393239;
   reg _393240_393240 ; 
   reg __393240_393240;
   reg _393241_393241 ; 
   reg __393241_393241;
   reg _393242_393242 ; 
   reg __393242_393242;
   reg _393243_393243 ; 
   reg __393243_393243;
   reg _393244_393244 ; 
   reg __393244_393244;
   reg _393245_393245 ; 
   reg __393245_393245;
   reg _393246_393246 ; 
   reg __393246_393246;
   reg _393247_393247 ; 
   reg __393247_393247;
   reg _393248_393248 ; 
   reg __393248_393248;
   reg _393249_393249 ; 
   reg __393249_393249;
   reg _393250_393250 ; 
   reg __393250_393250;
   reg _393251_393251 ; 
   reg __393251_393251;
   reg _393252_393252 ; 
   reg __393252_393252;
   reg _393253_393253 ; 
   reg __393253_393253;
   reg _393254_393254 ; 
   reg __393254_393254;
   reg _393255_393255 ; 
   reg __393255_393255;
   reg _393256_393256 ; 
   reg __393256_393256;
   reg _393257_393257 ; 
   reg __393257_393257;
   reg _393258_393258 ; 
   reg __393258_393258;
   reg _393259_393259 ; 
   reg __393259_393259;
   reg _393260_393260 ; 
   reg __393260_393260;
   reg _393261_393261 ; 
   reg __393261_393261;
   reg _393262_393262 ; 
   reg __393262_393262;
   reg _393263_393263 ; 
   reg __393263_393263;
   reg _393264_393264 ; 
   reg __393264_393264;
   reg _393265_393265 ; 
   reg __393265_393265;
   reg _393266_393266 ; 
   reg __393266_393266;
   reg _393267_393267 ; 
   reg __393267_393267;
   reg _393268_393268 ; 
   reg __393268_393268;
   reg _393269_393269 ; 
   reg __393269_393269;
   reg _393270_393270 ; 
   reg __393270_393270;
   reg _393271_393271 ; 
   reg __393271_393271;
   reg _393272_393272 ; 
   reg __393272_393272;
   reg _393273_393273 ; 
   reg __393273_393273;
   reg _393274_393274 ; 
   reg __393274_393274;
   reg _393275_393275 ; 
   reg __393275_393275;
   reg _393276_393276 ; 
   reg __393276_393276;
   reg _393277_393277 ; 
   reg __393277_393277;
   reg _393278_393278 ; 
   reg __393278_393278;
   reg _393279_393279 ; 
   reg __393279_393279;
   reg _393280_393280 ; 
   reg __393280_393280;
   reg _393281_393281 ; 
   reg __393281_393281;
   reg _393282_393282 ; 
   reg __393282_393282;
   reg _393283_393283 ; 
   reg __393283_393283;
   reg _393284_393284 ; 
   reg __393284_393284;
   reg _393285_393285 ; 
   reg __393285_393285;
   reg _393286_393286 ; 
   reg __393286_393286;
   reg _393287_393287 ; 
   reg __393287_393287;
   reg _393288_393288 ; 
   reg __393288_393288;
   reg _393289_393289 ; 
   reg __393289_393289;
   reg _393290_393290 ; 
   reg __393290_393290;
   reg _393291_393291 ; 
   reg __393291_393291;
   reg _393292_393292 ; 
   reg __393292_393292;
   reg _393293_393293 ; 
   reg __393293_393293;
   reg _393294_393294 ; 
   reg __393294_393294;
   reg _393295_393295 ; 
   reg __393295_393295;
   reg _393296_393296 ; 
   reg __393296_393296;
   reg _393297_393297 ; 
   reg __393297_393297;
   reg _393298_393298 ; 
   reg __393298_393298;
   reg _393299_393299 ; 
   reg __393299_393299;
   reg _393300_393300 ; 
   reg __393300_393300;
   reg _393301_393301 ; 
   reg __393301_393301;
   reg _393302_393302 ; 
   reg __393302_393302;
   reg _393303_393303 ; 
   reg __393303_393303;
   reg _393304_393304 ; 
   reg __393304_393304;
   reg _393305_393305 ; 
   reg __393305_393305;
   reg _393306_393306 ; 
   reg __393306_393306;
   reg _393307_393307 ; 
   reg __393307_393307;
   reg _393308_393308 ; 
   reg __393308_393308;
   reg _393309_393309 ; 
   reg __393309_393309;
   reg _393310_393310 ; 
   reg __393310_393310;
   reg _393311_393311 ; 
   reg __393311_393311;
   reg _393312_393312 ; 
   reg __393312_393312;
   reg _393313_393313 ; 
   reg __393313_393313;
   reg _393314_393314 ; 
   reg __393314_393314;
   reg _393315_393315 ; 
   reg __393315_393315;
   reg _393316_393316 ; 
   reg __393316_393316;
   reg _393317_393317 ; 
   reg __393317_393317;
   reg _393318_393318 ; 
   reg __393318_393318;
   reg _393319_393319 ; 
   reg __393319_393319;
   reg _393320_393320 ; 
   reg __393320_393320;
   reg _393321_393321 ; 
   reg __393321_393321;
   reg _393322_393322 ; 
   reg __393322_393322;
   reg _393323_393323 ; 
   reg __393323_393323;
   reg _393324_393324 ; 
   reg __393324_393324;
   reg _393325_393325 ; 
   reg __393325_393325;
   reg _393326_393326 ; 
   reg __393326_393326;
   reg _393327_393327 ; 
   reg __393327_393327;
   reg _393328_393328 ; 
   reg __393328_393328;
   reg _393329_393329 ; 
   reg __393329_393329;
   reg _393330_393330 ; 
   reg __393330_393330;
   reg _393331_393331 ; 
   reg __393331_393331;
   reg _393332_393332 ; 
   reg __393332_393332;
   reg _393333_393333 ; 
   reg __393333_393333;
   reg _393334_393334 ; 
   reg __393334_393334;
   reg _393335_393335 ; 
   reg __393335_393335;
   reg _393336_393336 ; 
   reg __393336_393336;
   reg _393337_393337 ; 
   reg __393337_393337;
   reg _393338_393338 ; 
   reg __393338_393338;
   reg _393339_393339 ; 
   reg __393339_393339;
   reg _393340_393340 ; 
   reg __393340_393340;
   reg _393341_393341 ; 
   reg __393341_393341;
   reg _393342_393342 ; 
   reg __393342_393342;
   reg _393343_393343 ; 
   reg __393343_393343;
   reg _393344_393344 ; 
   reg __393344_393344;
   reg _393345_393345 ; 
   reg __393345_393345;
   reg _393346_393346 ; 
   reg __393346_393346;
   reg _393347_393347 ; 
   reg __393347_393347;
   reg _393348_393348 ; 
   reg __393348_393348;
   reg _393349_393349 ; 
   reg __393349_393349;
   reg _393350_393350 ; 
   reg __393350_393350;
   reg _393351_393351 ; 
   reg __393351_393351;
   reg _393352_393352 ; 
   reg __393352_393352;
   reg _393353_393353 ; 
   reg __393353_393353;
   reg _393354_393354 ; 
   reg __393354_393354;
   reg _393355_393355 ; 
   reg __393355_393355;
   reg _393356_393356 ; 
   reg __393356_393356;
   reg _393357_393357 ; 
   reg __393357_393357;
   reg _393358_393358 ; 
   reg __393358_393358;
   reg _393359_393359 ; 
   reg __393359_393359;
   reg _393360_393360 ; 
   reg __393360_393360;
   reg _393361_393361 ; 
   reg __393361_393361;
   reg _393362_393362 ; 
   reg __393362_393362;
   reg _393363_393363 ; 
   reg __393363_393363;
   reg _393364_393364 ; 
   reg __393364_393364;
   reg _393365_393365 ; 
   reg __393365_393365;
   reg _393366_393366 ; 
   reg __393366_393366;
   reg _393367_393367 ; 
   reg __393367_393367;
   reg _393368_393368 ; 
   reg __393368_393368;
   reg _393369_393369 ; 
   reg __393369_393369;
   reg _393370_393370 ; 
   reg __393370_393370;
   reg _393371_393371 ; 
   reg __393371_393371;
   reg _393372_393372 ; 
   reg __393372_393372;
   reg _393373_393373 ; 
   reg __393373_393373;
   reg _393374_393374 ; 
   reg __393374_393374;
   reg _393375_393375 ; 
   reg __393375_393375;
   reg _393376_393376 ; 
   reg __393376_393376;
   reg _393377_393377 ; 
   reg __393377_393377;
   reg _393378_393378 ; 
   reg __393378_393378;
   reg _393379_393379 ; 
   reg __393379_393379;
   reg _393380_393380 ; 
   reg __393380_393380;
   reg _393381_393381 ; 
   reg __393381_393381;
   reg _393382_393382 ; 
   reg __393382_393382;
   reg _393383_393383 ; 
   reg __393383_393383;
   reg _393384_393384 ; 
   reg __393384_393384;
   reg _393385_393385 ; 
   reg __393385_393385;
   reg _393386_393386 ; 
   reg __393386_393386;
   reg _393387_393387 ; 
   reg __393387_393387;
   reg _393388_393388 ; 
   reg __393388_393388;
   reg _393389_393389 ; 
   reg __393389_393389;
   reg _393390_393390 ; 
   reg __393390_393390;
   reg _393391_393391 ; 
   reg __393391_393391;
   reg _393392_393392 ; 
   reg __393392_393392;
   reg _393393_393393 ; 
   reg __393393_393393;
   reg _393394_393394 ; 
   reg __393394_393394;
   reg _393395_393395 ; 
   reg __393395_393395;
   reg _393396_393396 ; 
   reg __393396_393396;
   reg _393397_393397 ; 
   reg __393397_393397;
   reg _393398_393398 ; 
   reg __393398_393398;
   reg _393399_393399 ; 
   reg __393399_393399;
   reg _393400_393400 ; 
   reg __393400_393400;
   reg _393401_393401 ; 
   reg __393401_393401;
   reg _393402_393402 ; 
   reg __393402_393402;
   reg _393403_393403 ; 
   reg __393403_393403;
   reg _393404_393404 ; 
   reg __393404_393404;
   reg _393405_393405 ; 
   reg __393405_393405;
   reg _393406_393406 ; 
   reg __393406_393406;
   reg _393407_393407 ; 
   reg __393407_393407;
   reg _393408_393408 ; 
   reg __393408_393408;
   reg _393409_393409 ; 
   reg __393409_393409;
   reg _393410_393410 ; 
   reg __393410_393410;
   reg _393411_393411 ; 
   reg __393411_393411;
   reg _393412_393412 ; 
   reg __393412_393412;
   reg _393413_393413 ; 
   reg __393413_393413;
   reg _393414_393414 ; 
   reg __393414_393414;
   reg _393415_393415 ; 
   reg __393415_393415;
   reg _393416_393416 ; 
   reg __393416_393416;
   reg _393417_393417 ; 
   reg __393417_393417;
   reg _393418_393418 ; 
   reg __393418_393418;
   reg _393419_393419 ; 
   reg __393419_393419;
   reg _393420_393420 ; 
   reg __393420_393420;
   reg _393421_393421 ; 
   reg __393421_393421;
   reg _393422_393422 ; 
   reg __393422_393422;
   reg _393423_393423 ; 
   reg __393423_393423;
   reg _393424_393424 ; 
   reg __393424_393424;
   reg _393425_393425 ; 
   reg __393425_393425;
   reg _393426_393426 ; 
   reg __393426_393426;
   reg _393427_393427 ; 
   reg __393427_393427;
   reg _393428_393428 ; 
   reg __393428_393428;
   reg _393429_393429 ; 
   reg __393429_393429;
   reg _393430_393430 ; 
   reg __393430_393430;
   reg _393431_393431 ; 
   reg __393431_393431;
   reg _393432_393432 ; 
   reg __393432_393432;
   reg _393433_393433 ; 
   reg __393433_393433;
   reg _393434_393434 ; 
   reg __393434_393434;
   reg _393435_393435 ; 
   reg __393435_393435;
   reg _393436_393436 ; 
   reg __393436_393436;
   reg _393437_393437 ; 
   reg __393437_393437;
   reg _393438_393438 ; 
   reg __393438_393438;
   reg _393439_393439 ; 
   reg __393439_393439;
   reg _393440_393440 ; 
   reg __393440_393440;
   reg _393441_393441 ; 
   reg __393441_393441;
   reg _393442_393442 ; 
   reg __393442_393442;
   reg _393443_393443 ; 
   reg __393443_393443;
   reg _393444_393444 ; 
   reg __393444_393444;
   reg _393445_393445 ; 
   reg __393445_393445;
   reg _393446_393446 ; 
   reg __393446_393446;
   reg _393447_393447 ; 
   reg __393447_393447;
   reg _393448_393448 ; 
   reg __393448_393448;
   reg _393449_393449 ; 
   reg __393449_393449;
   reg _393450_393450 ; 
   reg __393450_393450;
   reg _393451_393451 ; 
   reg __393451_393451;
   reg _393452_393452 ; 
   reg __393452_393452;
   reg _393453_393453 ; 
   reg __393453_393453;
   reg _393454_393454 ; 
   reg __393454_393454;
   reg _393455_393455 ; 
   reg __393455_393455;
   reg _393456_393456 ; 
   reg __393456_393456;
   reg _393457_393457 ; 
   reg __393457_393457;
   reg _393458_393458 ; 
   reg __393458_393458;
   reg _393459_393459 ; 
   reg __393459_393459;
   reg _393460_393460 ; 
   reg __393460_393460;
   reg _393461_393461 ; 
   reg __393461_393461;
   reg _393462_393462 ; 
   reg __393462_393462;
   reg _393463_393463 ; 
   reg __393463_393463;
   reg _393464_393464 ; 
   reg __393464_393464;
   reg _393465_393465 ; 
   reg __393465_393465;
   reg _393466_393466 ; 
   reg __393466_393466;
   reg _393467_393467 ; 
   reg __393467_393467;
   reg _393468_393468 ; 
   reg __393468_393468;
   reg _393469_393469 ; 
   reg __393469_393469;
   reg _393470_393470 ; 
   reg __393470_393470;
   reg _393471_393471 ; 
   reg __393471_393471;
   reg _393472_393472 ; 
   reg __393472_393472;
   reg _393473_393473 ; 
   reg __393473_393473;
   reg _393474_393474 ; 
   reg __393474_393474;
   reg _393475_393475 ; 
   reg __393475_393475;
   reg _393476_393476 ; 
   reg __393476_393476;
   reg _393477_393477 ; 
   reg __393477_393477;
   reg _393478_393478 ; 
   reg __393478_393478;
   reg _393479_393479 ; 
   reg __393479_393479;
   reg _393480_393480 ; 
   reg __393480_393480;
   reg _393481_393481 ; 
   reg __393481_393481;
   reg _393482_393482 ; 
   reg __393482_393482;
   reg _393483_393483 ; 
   reg __393483_393483;
   reg _393484_393484 ; 
   reg __393484_393484;
   reg _393485_393485 ; 
   reg __393485_393485;
   reg _393486_393486 ; 
   reg __393486_393486;
   reg _393487_393487 ; 
   reg __393487_393487;
   reg _393488_393488 ; 
   reg __393488_393488;
   reg _393489_393489 ; 
   reg __393489_393489;
   reg _393490_393490 ; 
   reg __393490_393490;
   reg _393491_393491 ; 
   reg __393491_393491;
   reg _393492_393492 ; 
   reg __393492_393492;
   reg _393493_393493 ; 
   reg __393493_393493;
   reg _393494_393494 ; 
   reg __393494_393494;
   reg _393495_393495 ; 
   reg __393495_393495;
   reg _393496_393496 ; 
   reg __393496_393496;
   reg _393497_393497 ; 
   reg __393497_393497;
   reg _393498_393498 ; 
   reg __393498_393498;
   reg _393499_393499 ; 
   reg __393499_393499;
   reg _393500_393500 ; 
   reg __393500_393500;
   reg _393501_393501 ; 
   reg __393501_393501;
   reg _393502_393502 ; 
   reg __393502_393502;
   reg _393503_393503 ; 
   reg __393503_393503;
   reg _393504_393504 ; 
   reg __393504_393504;
   reg _393505_393505 ; 
   reg __393505_393505;
   reg _393506_393506 ; 
   reg __393506_393506;
   reg _393507_393507 ; 
   reg __393507_393507;
   reg _393508_393508 ; 
   reg __393508_393508;
   reg _393509_393509 ; 
   reg __393509_393509;
   reg _393510_393510 ; 
   reg __393510_393510;
   reg _393511_393511 ; 
   reg __393511_393511;
   reg _393512_393512 ; 
   reg __393512_393512;
   reg _393513_393513 ; 
   reg __393513_393513;
   reg _393514_393514 ; 
   reg __393514_393514;
   reg _393515_393515 ; 
   reg __393515_393515;
   reg _393516_393516 ; 
   reg __393516_393516;
   reg _393517_393517 ; 
   reg __393517_393517;
   reg _393518_393518 ; 
   reg __393518_393518;
   reg _393519_393519 ; 
   reg __393519_393519;
   reg _393520_393520 ; 
   reg __393520_393520;
   reg _393521_393521 ; 
   reg __393521_393521;
   reg _393522_393522 ; 
   reg __393522_393522;
   reg _393523_393523 ; 
   reg __393523_393523;
   reg _393524_393524 ; 
   reg __393524_393524;
   reg _393525_393525 ; 
   reg __393525_393525;
   reg _393526_393526 ; 
   reg __393526_393526;
   reg _393527_393527 ; 
   reg __393527_393527;
   reg _393528_393528 ; 
   reg __393528_393528;
   reg _393529_393529 ; 
   reg __393529_393529;
   reg _393530_393530 ; 
   reg __393530_393530;
   reg _393531_393531 ; 
   reg __393531_393531;
   reg _393532_393532 ; 
   reg __393532_393532;
   reg _393533_393533 ; 
   reg __393533_393533;
   reg _393534_393534 ; 
   reg __393534_393534;
   reg _393535_393535 ; 
   reg __393535_393535;
   reg _393536_393536 ; 
   reg __393536_393536;
   reg _393537_393537 ; 
   reg __393537_393537;
   reg _393538_393538 ; 
   reg __393538_393538;
   reg _393539_393539 ; 
   reg __393539_393539;
   reg _393540_393540 ; 
   reg __393540_393540;
   reg _393541_393541 ; 
   reg __393541_393541;
   reg _393542_393542 ; 
   reg __393542_393542;
   reg _393543_393543 ; 
   reg __393543_393543;
   reg _393544_393544 ; 
   reg __393544_393544;
   reg _393545_393545 ; 
   reg __393545_393545;
   reg _393546_393546 ; 
   reg __393546_393546;
   reg _393547_393547 ; 
   reg __393547_393547;
   reg _393548_393548 ; 
   reg __393548_393548;
   reg _393549_393549 ; 
   reg __393549_393549;
   reg _393550_393550 ; 
   reg __393550_393550;
   reg _393551_393551 ; 
   reg __393551_393551;
   reg _393552_393552 ; 
   reg __393552_393552;
   reg _393553_393553 ; 
   reg __393553_393553;
   reg _393554_393554 ; 
   reg __393554_393554;
   reg _393555_393555 ; 
   reg __393555_393555;
   reg _393556_393556 ; 
   reg __393556_393556;
   reg _393557_393557 ; 
   reg __393557_393557;
   reg _393558_393558 ; 
   reg __393558_393558;
   reg _393559_393559 ; 
   reg __393559_393559;
   reg _393560_393560 ; 
   reg __393560_393560;
   reg _393561_393561 ; 
   reg __393561_393561;
   reg _393562_393562 ; 
   reg __393562_393562;
   reg _393563_393563 ; 
   reg __393563_393563;
   reg _393564_393564 ; 
   reg __393564_393564;
   reg _393565_393565 ; 
   reg __393565_393565;
   reg _393566_393566 ; 
   reg __393566_393566;
   reg _393567_393567 ; 
   reg __393567_393567;
   reg _393568_393568 ; 
   reg __393568_393568;
   reg _393569_393569 ; 
   reg __393569_393569;
   reg _393570_393570 ; 
   reg __393570_393570;
   reg _393571_393571 ; 
   reg __393571_393571;
   reg _393572_393572 ; 
   reg __393572_393572;
   reg _393573_393573 ; 
   reg __393573_393573;
   reg _393574_393574 ; 
   reg __393574_393574;
   reg _393575_393575 ; 
   reg __393575_393575;
   reg _393576_393576 ; 
   reg __393576_393576;
   reg _393577_393577 ; 
   reg __393577_393577;
   reg _393578_393578 ; 
   reg __393578_393578;
   reg _393579_393579 ; 
   reg __393579_393579;
   reg _393580_393580 ; 
   reg __393580_393580;
   reg _393581_393581 ; 
   reg __393581_393581;
   reg _393582_393582 ; 
   reg __393582_393582;
   reg _393583_393583 ; 
   reg __393583_393583;
   reg _393584_393584 ; 
   reg __393584_393584;
   reg _393585_393585 ; 
   reg __393585_393585;
   reg _393586_393586 ; 
   reg __393586_393586;
   reg _393587_393587 ; 
   reg __393587_393587;
   reg _393588_393588 ; 
   reg __393588_393588;
   reg _393589_393589 ; 
   reg __393589_393589;
   reg _393590_393590 ; 
   reg __393590_393590;
   reg _393591_393591 ; 
   reg __393591_393591;
   reg _393592_393592 ; 
   reg __393592_393592;
   reg _393593_393593 ; 
   reg __393593_393593;
   reg _393594_393594 ; 
   reg __393594_393594;
   reg _393595_393595 ; 
   reg __393595_393595;
   reg _393596_393596 ; 
   reg __393596_393596;
   reg _393597_393597 ; 
   reg __393597_393597;
   reg _393598_393598 ; 
   reg __393598_393598;
   reg _393599_393599 ; 
   reg __393599_393599;
   reg _393600_393600 ; 
   reg __393600_393600;
   reg _393601_393601 ; 
   reg __393601_393601;
   reg _393602_393602 ; 
   reg __393602_393602;
   reg _393603_393603 ; 
   reg __393603_393603;
   reg _393604_393604 ; 
   reg __393604_393604;
   reg _393605_393605 ; 
   reg __393605_393605;
   reg _393606_393606 ; 
   reg __393606_393606;
   reg _393607_393607 ; 
   reg __393607_393607;
   reg _393608_393608 ; 
   reg __393608_393608;
   reg _393609_393609 ; 
   reg __393609_393609;
   reg _393610_393610 ; 
   reg __393610_393610;
   reg _393611_393611 ; 
   reg __393611_393611;
   reg _393612_393612 ; 
   reg __393612_393612;
   reg _393613_393613 ; 
   reg __393613_393613;
   reg _393614_393614 ; 
   reg __393614_393614;
   reg _393615_393615 ; 
   reg __393615_393615;
   reg _393616_393616 ; 
   reg __393616_393616;
   reg _393617_393617 ; 
   reg __393617_393617;
   reg _393618_393618 ; 
   reg __393618_393618;
   reg _393619_393619 ; 
   reg __393619_393619;
   reg _393620_393620 ; 
   reg __393620_393620;
   reg _393621_393621 ; 
   reg __393621_393621;
   reg _393622_393622 ; 
   reg __393622_393622;
   reg _393623_393623 ; 
   reg __393623_393623;
   reg _393624_393624 ; 
   reg __393624_393624;
   reg _393625_393625 ; 
   reg __393625_393625;
   reg _393626_393626 ; 
   reg __393626_393626;
   reg _393627_393627 ; 
   reg __393627_393627;
   reg _393628_393628 ; 
   reg __393628_393628;
   reg _393629_393629 ; 
   reg __393629_393629;
   reg _393630_393630 ; 
   reg __393630_393630;
   reg _393631_393631 ; 
   reg __393631_393631;
   reg _393632_393632 ; 
   reg __393632_393632;
   reg _393633_393633 ; 
   reg __393633_393633;
   reg _393634_393634 ; 
   reg __393634_393634;
   reg _393635_393635 ; 
   reg __393635_393635;
   reg _393636_393636 ; 
   reg __393636_393636;
   reg _393637_393637 ; 
   reg __393637_393637;
   reg _393638_393638 ; 
   reg __393638_393638;
   reg _393639_393639 ; 
   reg __393639_393639;
   reg _393640_393640 ; 
   reg __393640_393640;
   reg _393641_393641 ; 
   reg __393641_393641;
   reg _393642_393642 ; 
   reg __393642_393642;
   reg _393643_393643 ; 
   reg __393643_393643;
   reg _393644_393644 ; 
   reg __393644_393644;
   reg _393645_393645 ; 
   reg __393645_393645;
   reg _393646_393646 ; 
   reg __393646_393646;
   reg _393647_393647 ; 
   reg __393647_393647;
   reg _393648_393648 ; 
   reg __393648_393648;
   reg _393649_393649 ; 
   reg __393649_393649;
   reg _393650_393650 ; 
   reg __393650_393650;
   reg _393651_393651 ; 
   reg __393651_393651;
   reg _393652_393652 ; 
   reg __393652_393652;
   reg _393653_393653 ; 
   reg __393653_393653;
   reg _393654_393654 ; 
   reg __393654_393654;
   reg _393655_393655 ; 
   reg __393655_393655;
   reg _393656_393656 ; 
   reg __393656_393656;
   reg _393657_393657 ; 
   reg __393657_393657;
   reg _393658_393658 ; 
   reg __393658_393658;
   reg _393659_393659 ; 
   reg __393659_393659;
   reg _393660_393660 ; 
   reg __393660_393660;
   reg _393661_393661 ; 
   reg __393661_393661;
   reg _393662_393662 ; 
   reg __393662_393662;
   reg _393663_393663 ; 
   reg __393663_393663;
   reg _393664_393664 ; 
   reg __393664_393664;
   reg _393665_393665 ; 
   reg __393665_393665;
   reg _393666_393666 ; 
   reg __393666_393666;
   reg _393667_393667 ; 
   reg __393667_393667;
   reg _393668_393668 ; 
   reg __393668_393668;
   reg _393669_393669 ; 
   reg __393669_393669;
   reg _393670_393670 ; 
   reg __393670_393670;
   reg _393671_393671 ; 
   reg __393671_393671;
   reg _393672_393672 ; 
   reg __393672_393672;
   reg _393673_393673 ; 
   reg __393673_393673;
   reg _393674_393674 ; 
   reg __393674_393674;
   reg _393675_393675 ; 
   reg __393675_393675;
   reg _393676_393676 ; 
   reg __393676_393676;
   reg _393677_393677 ; 
   reg __393677_393677;
   reg _393678_393678 ; 
   reg __393678_393678;
   reg _393679_393679 ; 
   reg __393679_393679;
   reg _393680_393680 ; 
   reg __393680_393680;
   reg _393681_393681 ; 
   reg __393681_393681;
   reg _393682_393682 ; 
   reg __393682_393682;
   reg _393683_393683 ; 
   reg __393683_393683;
   reg _393684_393684 ; 
   reg __393684_393684;
   reg _393685_393685 ; 
   reg __393685_393685;
   reg _393686_393686 ; 
   reg __393686_393686;
   reg _393687_393687 ; 
   reg __393687_393687;
   reg _393688_393688 ; 
   reg __393688_393688;
   reg _393689_393689 ; 
   reg __393689_393689;
   reg _393690_393690 ; 
   reg __393690_393690;
   reg _393691_393691 ; 
   reg __393691_393691;
   reg _393692_393692 ; 
   reg __393692_393692;
   reg _393693_393693 ; 
   reg __393693_393693;
   reg _393694_393694 ; 
   reg __393694_393694;
   reg _393695_393695 ; 
   reg __393695_393695;
   reg _393696_393696 ; 
   reg __393696_393696;
   reg _393697_393697 ; 
   reg __393697_393697;
   reg _393698_393698 ; 
   reg __393698_393698;
   reg _393699_393699 ; 
   reg __393699_393699;
   reg _393700_393700 ; 
   reg __393700_393700;
   reg _393701_393701 ; 
   reg __393701_393701;
   reg _393702_393702 ; 
   reg __393702_393702;
   reg _393703_393703 ; 
   reg __393703_393703;
   reg _393704_393704 ; 
   reg __393704_393704;
   reg _393705_393705 ; 
   reg __393705_393705;
   reg _393706_393706 ; 
   reg __393706_393706;
   reg _393707_393707 ; 
   reg __393707_393707;
   reg _393708_393708 ; 
   reg __393708_393708;
   reg _393709_393709 ; 
   reg __393709_393709;
   reg _393710_393710 ; 
   reg __393710_393710;
   reg _393711_393711 ; 
   reg __393711_393711;
   reg _393712_393712 ; 
   reg __393712_393712;
   reg _393713_393713 ; 
   reg __393713_393713;
   reg _393714_393714 ; 
   reg __393714_393714;
   reg _393715_393715 ; 
   reg __393715_393715;
   reg _393716_393716 ; 
   reg __393716_393716;
   reg _393717_393717 ; 
   reg __393717_393717;
   reg _393718_393718 ; 
   reg __393718_393718;
   reg _393719_393719 ; 
   reg __393719_393719;
   reg _393720_393720 ; 
   reg __393720_393720;
   reg _393721_393721 ; 
   reg __393721_393721;
   reg _393722_393722 ; 
   reg __393722_393722;
   reg _393723_393723 ; 
   reg __393723_393723;
   reg _393724_393724 ; 
   reg __393724_393724;
   reg _393725_393725 ; 
   reg __393725_393725;
   reg _393726_393726 ; 
   reg __393726_393726;
   reg _393727_393727 ; 
   reg __393727_393727;
   reg _393728_393728 ; 
   reg __393728_393728;
   reg _393729_393729 ; 
   reg __393729_393729;
   reg _393730_393730 ; 
   reg __393730_393730;
   reg _393731_393731 ; 
   reg __393731_393731;
   reg _393732_393732 ; 
   reg __393732_393732;
   reg _393733_393733 ; 
   reg __393733_393733;
   reg _393734_393734 ; 
   reg __393734_393734;
   reg _393735_393735 ; 
   reg __393735_393735;
   reg _393736_393736 ; 
   reg __393736_393736;
   reg _393737_393737 ; 
   reg __393737_393737;
   reg _393738_393738 ; 
   reg __393738_393738;
   reg _393739_393739 ; 
   reg __393739_393739;
   reg _393740_393740 ; 
   reg __393740_393740;
   reg _393741_393741 ; 
   reg __393741_393741;
   reg _393742_393742 ; 
   reg __393742_393742;
   reg _393743_393743 ; 
   reg __393743_393743;
   reg _393744_393744 ; 
   reg __393744_393744;
   reg _393745_393745 ; 
   reg __393745_393745;
   reg _393746_393746 ; 
   reg __393746_393746;
   reg _393747_393747 ; 
   reg __393747_393747;
   reg _393748_393748 ; 
   reg __393748_393748;
   reg _393749_393749 ; 
   reg __393749_393749;
   reg _393750_393750 ; 
   reg __393750_393750;
   reg _393751_393751 ; 
   reg __393751_393751;
   reg _393752_393752 ; 
   reg __393752_393752;
   reg _393753_393753 ; 
   reg __393753_393753;
   reg _393754_393754 ; 
   reg __393754_393754;
   reg _393755_393755 ; 
   reg __393755_393755;
   reg _393756_393756 ; 
   reg __393756_393756;
   reg _393757_393757 ; 
   reg __393757_393757;
   reg _393758_393758 ; 
   reg __393758_393758;
   reg _393759_393759 ; 
   reg __393759_393759;
   reg _393760_393760 ; 
   reg __393760_393760;
   reg _393761_393761 ; 
   reg __393761_393761;
   reg _393762_393762 ; 
   reg __393762_393762;
   reg _393763_393763 ; 
   reg __393763_393763;
   reg _393764_393764 ; 
   reg __393764_393764;
   reg _393765_393765 ; 
   reg __393765_393765;
   reg _393766_393766 ; 
   reg __393766_393766;
   reg _393767_393767 ; 
   reg __393767_393767;
   reg _393768_393768 ; 
   reg __393768_393768;
   reg _393769_393769 ; 
   reg __393769_393769;
   reg _393770_393770 ; 
   reg __393770_393770;
   reg _393771_393771 ; 
   reg __393771_393771;
   reg _393772_393772 ; 
   reg __393772_393772;
   reg _393773_393773 ; 
   reg __393773_393773;
   reg _393774_393774 ; 
   reg __393774_393774;
   reg _393775_393775 ; 
   reg __393775_393775;
   reg _393776_393776 ; 
   reg __393776_393776;
   reg _393777_393777 ; 
   reg __393777_393777;
   reg _393778_393778 ; 
   reg __393778_393778;
   reg _393779_393779 ; 
   reg __393779_393779;
   reg _393780_393780 ; 
   reg __393780_393780;
   reg _393781_393781 ; 
   reg __393781_393781;
   reg _393782_393782 ; 
   reg __393782_393782;
   reg _393783_393783 ; 
   reg __393783_393783;
   reg _393784_393784 ; 
   reg __393784_393784;
   reg _393785_393785 ; 
   reg __393785_393785;
   reg _393786_393786 ; 
   reg __393786_393786;
   reg _393787_393787 ; 
   reg __393787_393787;
   reg _393788_393788 ; 
   reg __393788_393788;
   reg _393789_393789 ; 
   reg __393789_393789;
   reg _393790_393790 ; 
   reg __393790_393790;
   reg _393791_393791 ; 
   reg __393791_393791;
   reg _393792_393792 ; 
   reg __393792_393792;
   reg _393793_393793 ; 
   reg __393793_393793;
   reg _393794_393794 ; 
   reg __393794_393794;
   reg _393795_393795 ; 
   reg __393795_393795;
   reg _393796_393796 ; 
   reg __393796_393796;
   reg _393797_393797 ; 
   reg __393797_393797;
   reg _393798_393798 ; 
   reg __393798_393798;
   reg _393799_393799 ; 
   reg __393799_393799;
   reg _393800_393800 ; 
   reg __393800_393800;
   reg _393801_393801 ; 
   reg __393801_393801;
   reg _393802_393802 ; 
   reg __393802_393802;
   reg _393803_393803 ; 
   reg __393803_393803;
   reg _393804_393804 ; 
   reg __393804_393804;
   reg _393805_393805 ; 
   reg __393805_393805;
   reg _393806_393806 ; 
   reg __393806_393806;
   reg _393807_393807 ; 
   reg __393807_393807;
   reg _393808_393808 ; 
   reg __393808_393808;
   reg _393809_393809 ; 
   reg __393809_393809;
   reg _393810_393810 ; 
   reg __393810_393810;
   reg _393811_393811 ; 
   reg __393811_393811;
   reg _393812_393812 ; 
   reg __393812_393812;
   reg _393813_393813 ; 
   reg __393813_393813;
   reg _393814_393814 ; 
   reg __393814_393814;
   reg _393815_393815 ; 
   reg __393815_393815;
   reg _393816_393816 ; 
   reg __393816_393816;
   reg _393817_393817 ; 
   reg __393817_393817;
   reg _393818_393818 ; 
   reg __393818_393818;
   reg _393819_393819 ; 
   reg __393819_393819;
   reg _393820_393820 ; 
   reg __393820_393820;
   reg _393821_393821 ; 
   reg __393821_393821;
   reg _393822_393822 ; 
   reg __393822_393822;
   reg _393823_393823 ; 
   reg __393823_393823;
   reg _393824_393824 ; 
   reg __393824_393824;
   reg _393825_393825 ; 
   reg __393825_393825;
   reg _393826_393826 ; 
   reg __393826_393826;
   reg _393827_393827 ; 
   reg __393827_393827;
   reg _393828_393828 ; 
   reg __393828_393828;
   reg _393829_393829 ; 
   reg __393829_393829;
   reg _393830_393830 ; 
   reg __393830_393830;
   reg _393831_393831 ; 
   reg __393831_393831;
   reg _393832_393832 ; 
   reg __393832_393832;
   reg _393833_393833 ; 
   reg __393833_393833;
   reg _393834_393834 ; 
   reg __393834_393834;
   reg _393835_393835 ; 
   reg __393835_393835;
   reg _393836_393836 ; 
   reg __393836_393836;
   reg _393837_393837 ; 
   reg __393837_393837;
   reg _393838_393838 ; 
   reg __393838_393838;
   reg _393839_393839 ; 
   reg __393839_393839;
   reg _393840_393840 ; 
   reg __393840_393840;
   reg _393841_393841 ; 
   reg __393841_393841;
   reg _393842_393842 ; 
   reg __393842_393842;
   reg _393843_393843 ; 
   reg __393843_393843;
   reg _393844_393844 ; 
   reg __393844_393844;
   reg _393845_393845 ; 
   reg __393845_393845;
   reg _393846_393846 ; 
   reg __393846_393846;
   reg _393847_393847 ; 
   reg __393847_393847;
   reg _393848_393848 ; 
   reg __393848_393848;
   reg _393849_393849 ; 
   reg __393849_393849;
   reg _393850_393850 ; 
   reg __393850_393850;
   reg _393851_393851 ; 
   reg __393851_393851;
   reg _393852_393852 ; 
   reg __393852_393852;
   reg _393853_393853 ; 
   reg __393853_393853;
   reg _393854_393854 ; 
   reg __393854_393854;
   reg _393855_393855 ; 
   reg __393855_393855;
   reg _393856_393856 ; 
   reg __393856_393856;
   reg _393857_393857 ; 
   reg __393857_393857;
   reg _393858_393858 ; 
   reg __393858_393858;
   reg _393859_393859 ; 
   reg __393859_393859;
   reg _393860_393860 ; 
   reg __393860_393860;
   reg _393861_393861 ; 
   reg __393861_393861;
   reg _393862_393862 ; 
   reg __393862_393862;
   reg _393863_393863 ; 
   reg __393863_393863;
   reg _393864_393864 ; 
   reg __393864_393864;
   reg _393865_393865 ; 
   reg __393865_393865;
   reg _393866_393866 ; 
   reg __393866_393866;
   reg _393867_393867 ; 
   reg __393867_393867;
   reg _393868_393868 ; 
   reg __393868_393868;
   reg _393869_393869 ; 
   reg __393869_393869;
   reg _393870_393870 ; 
   reg __393870_393870;
   reg _393871_393871 ; 
   reg __393871_393871;
   reg _393872_393872 ; 
   reg __393872_393872;
   reg _393873_393873 ; 
   reg __393873_393873;
   reg _393874_393874 ; 
   reg __393874_393874;
   reg _393875_393875 ; 
   reg __393875_393875;
   reg _393876_393876 ; 
   reg __393876_393876;
   reg _393877_393877 ; 
   reg __393877_393877;
   reg _393878_393878 ; 
   reg __393878_393878;
   reg _393879_393879 ; 
   reg __393879_393879;
   reg _393880_393880 ; 
   reg __393880_393880;
   reg _393881_393881 ; 
   reg __393881_393881;
   reg _393882_393882 ; 
   reg __393882_393882;
   reg _393883_393883 ; 
   reg __393883_393883;
   reg _393884_393884 ; 
   reg __393884_393884;
   reg _393885_393885 ; 
   reg __393885_393885;
   reg _393886_393886 ; 
   reg __393886_393886;
   reg _393887_393887 ; 
   reg __393887_393887;
   reg _393888_393888 ; 
   reg __393888_393888;
   reg _393889_393889 ; 
   reg __393889_393889;
   reg _393890_393890 ; 
   reg __393890_393890;
   reg _393891_393891 ; 
   reg __393891_393891;
   reg _393892_393892 ; 
   reg __393892_393892;
   reg _393893_393893 ; 
   reg __393893_393893;
   reg _393894_393894 ; 
   reg __393894_393894;
   reg _393895_393895 ; 
   reg __393895_393895;
   reg _393896_393896 ; 
   reg __393896_393896;
   reg _393897_393897 ; 
   reg __393897_393897;
   reg _393898_393898 ; 
   reg __393898_393898;
   reg _393899_393899 ; 
   reg __393899_393899;
   reg _393900_393900 ; 
   reg __393900_393900;
   reg _393901_393901 ; 
   reg __393901_393901;
   reg _393902_393902 ; 
   reg __393902_393902;
   reg _393903_393903 ; 
   reg __393903_393903;
   reg _393904_393904 ; 
   reg __393904_393904;
   reg _393905_393905 ; 
   reg __393905_393905;
   reg _393906_393906 ; 
   reg __393906_393906;
   reg _393907_393907 ; 
   reg __393907_393907;
   reg _393908_393908 ; 
   reg __393908_393908;
   reg _393909_393909 ; 
   reg __393909_393909;
   reg _393910_393910 ; 
   reg __393910_393910;
   reg _393911_393911 ; 
   reg __393911_393911;
   reg _393912_393912 ; 
   reg __393912_393912;
   reg _393913_393913 ; 
   reg __393913_393913;
   reg _393914_393914 ; 
   reg __393914_393914;
   reg _393915_393915 ; 
   reg __393915_393915;
   reg _393916_393916 ; 
   reg __393916_393916;
   reg _393917_393917 ; 
   reg __393917_393917;
   reg _393918_393918 ; 
   reg __393918_393918;
   reg _393919_393919 ; 
   reg __393919_393919;
   reg _393920_393920 ; 
   reg __393920_393920;
   reg _393921_393921 ; 
   reg __393921_393921;
   reg _393922_393922 ; 
   reg __393922_393922;
   reg _393923_393923 ; 
   reg __393923_393923;
   reg _393924_393924 ; 
   reg __393924_393924;
   reg _393925_393925 ; 
   reg __393925_393925;
   reg _393926_393926 ; 
   reg __393926_393926;
   reg _393927_393927 ; 
   reg __393927_393927;
   reg _393928_393928 ; 
   reg __393928_393928;
   reg _393929_393929 ; 
   reg __393929_393929;
   reg _393930_393930 ; 
   reg __393930_393930;
   reg _393931_393931 ; 
   reg __393931_393931;
   reg _393932_393932 ; 
   reg __393932_393932;
   reg _393933_393933 ; 
   reg __393933_393933;
   reg _393934_393934 ; 
   reg __393934_393934;
   reg _393935_393935 ; 
   reg __393935_393935;
   reg _393936_393936 ; 
   reg __393936_393936;
   reg _393937_393937 ; 
   reg __393937_393937;
   reg _393938_393938 ; 
   reg __393938_393938;
   reg _393939_393939 ; 
   reg __393939_393939;
   reg _393940_393940 ; 
   reg __393940_393940;
   reg _393941_393941 ; 
   reg __393941_393941;
   reg _393942_393942 ; 
   reg __393942_393942;
   reg _393943_393943 ; 
   reg __393943_393943;
   reg _393944_393944 ; 
   reg __393944_393944;
   reg _393945_393945 ; 
   reg __393945_393945;
   reg _393946_393946 ; 
   reg __393946_393946;
   reg _393947_393947 ; 
   reg __393947_393947;
   reg _393948_393948 ; 
   reg __393948_393948;
   reg _393949_393949 ; 
   reg __393949_393949;
   reg _393950_393950 ; 
   reg __393950_393950;
   reg _393951_393951 ; 
   reg __393951_393951;
   reg _393952_393952 ; 
   reg __393952_393952;
   reg _393953_393953 ; 
   reg __393953_393953;
   reg _393954_393954 ; 
   reg __393954_393954;
   reg _393955_393955 ; 
   reg __393955_393955;
   reg _393956_393956 ; 
   reg __393956_393956;
   reg _393957_393957 ; 
   reg __393957_393957;
   reg _393958_393958 ; 
   reg __393958_393958;
   reg _393959_393959 ; 
   reg __393959_393959;
   reg _393960_393960 ; 
   reg __393960_393960;
   reg _393961_393961 ; 
   reg __393961_393961;
   reg _393962_393962 ; 
   reg __393962_393962;
   reg _393963_393963 ; 
   reg __393963_393963;
   reg _393964_393964 ; 
   reg __393964_393964;
   reg _393965_393965 ; 
   reg __393965_393965;
   reg _393966_393966 ; 
   reg __393966_393966;
   reg _393967_393967 ; 
   reg __393967_393967;
   reg _393968_393968 ; 
   reg __393968_393968;
   reg _393969_393969 ; 
   reg __393969_393969;
   reg _393970_393970 ; 
   reg __393970_393970;
   reg _393971_393971 ; 
   reg __393971_393971;
   reg _393972_393972 ; 
   reg __393972_393972;
   reg _393973_393973 ; 
   reg __393973_393973;
   reg _393974_393974 ; 
   reg __393974_393974;
   reg _393975_393975 ; 
   reg __393975_393975;
   reg _393976_393976 ; 
   reg __393976_393976;
   reg _393977_393977 ; 
   reg __393977_393977;
   reg _393978_393978 ; 
   reg __393978_393978;
   reg _393979_393979 ; 
   reg __393979_393979;
   reg _393980_393980 ; 
   reg __393980_393980;
   reg _393981_393981 ; 
   reg __393981_393981;
   reg _393982_393982 ; 
   reg __393982_393982;
   reg _393983_393983 ; 
   reg __393983_393983;
   reg _393984_393984 ; 
   reg __393984_393984;
   reg _393985_393985 ; 
   reg __393985_393985;
   reg _393986_393986 ; 
   reg __393986_393986;
   reg _393987_393987 ; 
   reg __393987_393987;
   reg _393988_393988 ; 
   reg __393988_393988;
   reg _393989_393989 ; 
   reg __393989_393989;
   reg _393990_393990 ; 
   reg __393990_393990;
   reg _393991_393991 ; 
   reg __393991_393991;
   reg _393992_393992 ; 
   reg __393992_393992;
   reg _393993_393993 ; 
   reg __393993_393993;
   reg _393994_393994 ; 
   reg __393994_393994;
   reg _393995_393995 ; 
   reg __393995_393995;
   reg _393996_393996 ; 
   reg __393996_393996;
   reg _393997_393997 ; 
   reg __393997_393997;
   reg _393998_393998 ; 
   reg __393998_393998;
   reg _393999_393999 ; 
   reg __393999_393999;
   reg _394000_394000 ; 
   reg __394000_394000;
   reg _394001_394001 ; 
   reg __394001_394001;
   reg _394002_394002 ; 
   reg __394002_394002;
   reg _394003_394003 ; 
   reg __394003_394003;
   reg _394004_394004 ; 
   reg __394004_394004;
   reg _394005_394005 ; 
   reg __394005_394005;
   reg _394006_394006 ; 
   reg __394006_394006;
   reg _394007_394007 ; 
   reg __394007_394007;
   reg _394008_394008 ; 
   reg __394008_394008;
   reg _394009_394009 ; 
   reg __394009_394009;
   reg _394010_394010 ; 
   reg __394010_394010;
   reg _394011_394011 ; 
   reg __394011_394011;
   reg _394012_394012 ; 
   reg __394012_394012;
   reg _394013_394013 ; 
   reg __394013_394013;
   reg _394014_394014 ; 
   reg __394014_394014;
   reg _394015_394015 ; 
   reg __394015_394015;
   reg _394016_394016 ; 
   reg __394016_394016;
   reg _394017_394017 ; 
   reg __394017_394017;
   reg _394018_394018 ; 
   reg __394018_394018;
   reg _394019_394019 ; 
   reg __394019_394019;
   reg _394020_394020 ; 
   reg __394020_394020;
   reg _394021_394021 ; 
   reg __394021_394021;
   reg _394022_394022 ; 
   reg __394022_394022;
   reg _394023_394023 ; 
   reg __394023_394023;
   reg _394024_394024 ; 
   reg __394024_394024;
   reg _394025_394025 ; 
   reg __394025_394025;
   reg _394026_394026 ; 
   reg __394026_394026;
   reg _394027_394027 ; 
   reg __394027_394027;
   reg _394028_394028 ; 
   reg __394028_394028;
   reg _394029_394029 ; 
   reg __394029_394029;
   reg _394030_394030 ; 
   reg __394030_394030;
   reg _394031_394031 ; 
   reg __394031_394031;
   reg _394032_394032 ; 
   reg __394032_394032;
   reg _394033_394033 ; 
   reg __394033_394033;
   reg _394034_394034 ; 
   reg __394034_394034;
   reg _394035_394035 ; 
   reg __394035_394035;
   reg _394036_394036 ; 
   reg __394036_394036;
   reg _394037_394037 ; 
   reg __394037_394037;
   reg _394038_394038 ; 
   reg __394038_394038;
   reg _394039_394039 ; 
   reg __394039_394039;
   reg _394040_394040 ; 
   reg __394040_394040;
   reg _394041_394041 ; 
   reg __394041_394041;
   reg _394042_394042 ; 
   reg __394042_394042;
   reg _394043_394043 ; 
   reg __394043_394043;
   reg _394044_394044 ; 
   reg __394044_394044;
   reg _394045_394045 ; 
   reg __394045_394045;
   reg _394046_394046 ; 
   reg __394046_394046;
   reg _394047_394047 ; 
   reg __394047_394047;
   reg _394048_394048 ; 
   reg __394048_394048;
   reg _394049_394049 ; 
   reg __394049_394049;
   reg _394050_394050 ; 
   reg __394050_394050;
   reg _394051_394051 ; 
   reg __394051_394051;
   reg _394052_394052 ; 
   reg __394052_394052;
   reg _394053_394053 ; 
   reg __394053_394053;
   reg _394054_394054 ; 
   reg __394054_394054;
   reg _394055_394055 ; 
   reg __394055_394055;
   reg _394056_394056 ; 
   reg __394056_394056;
   reg _394057_394057 ; 
   reg __394057_394057;
   reg _394058_394058 ; 
   reg __394058_394058;
   reg _394059_394059 ; 
   reg __394059_394059;
   reg _394060_394060 ; 
   reg __394060_394060;
   reg _394061_394061 ; 
   reg __394061_394061;
   reg _394062_394062 ; 
   reg __394062_394062;
   reg _394063_394063 ; 
   reg __394063_394063;
   reg _394064_394064 ; 
   reg __394064_394064;
   reg _394065_394065 ; 
   reg __394065_394065;
   reg _394066_394066 ; 
   reg __394066_394066;
   reg _394067_394067 ; 
   reg __394067_394067;
   reg _394068_394068 ; 
   reg __394068_394068;
   reg _394069_394069 ; 
   reg __394069_394069;
   reg _394070_394070 ; 
   reg __394070_394070;
   reg _394071_394071 ; 
   reg __394071_394071;
   reg _394072_394072 ; 
   reg __394072_394072;
   reg _394073_394073 ; 
   reg __394073_394073;
   reg _394074_394074 ; 
   reg __394074_394074;
   reg _394075_394075 ; 
   reg __394075_394075;
   reg _394076_394076 ; 
   reg __394076_394076;
   reg _394077_394077 ; 
   reg __394077_394077;
   reg _394078_394078 ; 
   reg __394078_394078;
   reg _394079_394079 ; 
   reg __394079_394079;
   reg _394080_394080 ; 
   reg __394080_394080;
   reg _394081_394081 ; 
   reg __394081_394081;
   reg _394082_394082 ; 
   reg __394082_394082;
   reg _394083_394083 ; 
   reg __394083_394083;
   reg _394084_394084 ; 
   reg __394084_394084;
   reg _394085_394085 ; 
   reg __394085_394085;
   reg _394086_394086 ; 
   reg __394086_394086;
   reg _394087_394087 ; 
   reg __394087_394087;
   reg _394088_394088 ; 
   reg __394088_394088;
   reg _394089_394089 ; 
   reg __394089_394089;
   reg _394090_394090 ; 
   reg __394090_394090;
   reg _394091_394091 ; 
   reg __394091_394091;
   reg _394092_394092 ; 
   reg __394092_394092;
   reg _394093_394093 ; 
   reg __394093_394093;
   reg _394094_394094 ; 
   reg __394094_394094;
   reg _394095_394095 ; 
   reg __394095_394095;
   reg _394096_394096 ; 
   reg __394096_394096;
   reg _394097_394097 ; 
   reg __394097_394097;
   reg _394098_394098 ; 
   reg __394098_394098;
   reg _394099_394099 ; 
   reg __394099_394099;
   reg _394100_394100 ; 
   reg __394100_394100;
   reg _394101_394101 ; 
   reg __394101_394101;
   reg _394102_394102 ; 
   reg __394102_394102;
   reg _394103_394103 ; 
   reg __394103_394103;
   reg _394104_394104 ; 
   reg __394104_394104;
   reg _394105_394105 ; 
   reg __394105_394105;
   reg _394106_394106 ; 
   reg __394106_394106;
   reg _394107_394107 ; 
   reg __394107_394107;
   reg _394108_394108 ; 
   reg __394108_394108;
   reg _394109_394109 ; 
   reg __394109_394109;
   reg _394110_394110 ; 
   reg __394110_394110;
   reg _394111_394111 ; 
   reg __394111_394111;
   reg _394112_394112 ; 
   reg __394112_394112;
   reg _394113_394113 ; 
   reg __394113_394113;
   reg _394114_394114 ; 
   reg __394114_394114;
   reg _394115_394115 ; 
   reg __394115_394115;
   reg _394116_394116 ; 
   reg __394116_394116;
   reg _394117_394117 ; 
   reg __394117_394117;
   reg _394118_394118 ; 
   reg __394118_394118;
   reg _394119_394119 ; 
   reg __394119_394119;
   reg _394120_394120 ; 
   reg __394120_394120;
   reg _394121_394121 ; 
   reg __394121_394121;
   reg _394122_394122 ; 
   reg __394122_394122;
   reg _394123_394123 ; 
   reg __394123_394123;
   reg _394124_394124 ; 
   reg __394124_394124;
   reg _394125_394125 ; 
   reg __394125_394125;
   reg _394126_394126 ; 
   reg __394126_394126;
   reg _394127_394127 ; 
   reg __394127_394127;
   reg _394128_394128 ; 
   reg __394128_394128;
   reg _394129_394129 ; 
   reg __394129_394129;
   reg _394130_394130 ; 
   reg __394130_394130;
   reg _394131_394131 ; 
   reg __394131_394131;
   reg _394132_394132 ; 
   reg __394132_394132;
   reg _394133_394133 ; 
   reg __394133_394133;
   reg _394134_394134 ; 
   reg __394134_394134;
   reg _394135_394135 ; 
   reg __394135_394135;
   reg _394136_394136 ; 
   reg __394136_394136;
   reg _394137_394137 ; 
   reg __394137_394137;
   reg _394138_394138 ; 
   reg __394138_394138;
   reg _394139_394139 ; 
   reg __394139_394139;
   reg _394140_394140 ; 
   reg __394140_394140;
   reg _394141_394141 ; 
   reg __394141_394141;
   reg _394142_394142 ; 
   reg __394142_394142;
   reg _394143_394143 ; 
   reg __394143_394143;
   reg _394144_394144 ; 
   reg __394144_394144;
   reg _394145_394145 ; 
   reg __394145_394145;
   reg _394146_394146 ; 
   reg __394146_394146;
   reg _394147_394147 ; 
   reg __394147_394147;
   reg _394148_394148 ; 
   reg __394148_394148;
   reg _394149_394149 ; 
   reg __394149_394149;
   reg _394150_394150 ; 
   reg __394150_394150;
   reg _394151_394151 ; 
   reg __394151_394151;
   reg _394152_394152 ; 
   reg __394152_394152;
   reg _394153_394153 ; 
   reg __394153_394153;
   reg _394154_394154 ; 
   reg __394154_394154;
   reg _394155_394155 ; 
   reg __394155_394155;
   reg _394156_394156 ; 
   reg __394156_394156;
   reg _394157_394157 ; 
   reg __394157_394157;
   reg _394158_394158 ; 
   reg __394158_394158;
   reg _394159_394159 ; 
   reg __394159_394159;
   reg _394160_394160 ; 
   reg __394160_394160;
   reg _394161_394161 ; 
   reg __394161_394161;
   reg _394162_394162 ; 
   reg __394162_394162;
   reg _394163_394163 ; 
   reg __394163_394163;
   reg _394164_394164 ; 
   reg __394164_394164;
   reg _394165_394165 ; 
   reg __394165_394165;
   reg _394166_394166 ; 
   reg __394166_394166;
   reg _394167_394167 ; 
   reg __394167_394167;
   reg _394168_394168 ; 
   reg __394168_394168;
   reg _394169_394169 ; 
   reg __394169_394169;
   reg _394170_394170 ; 
   reg __394170_394170;
   reg _394171_394171 ; 
   reg __394171_394171;
   reg _394172_394172 ; 
   reg __394172_394172;
   reg _394173_394173 ; 
   reg __394173_394173;
   reg _394174_394174 ; 
   reg __394174_394174;
   reg _394175_394175 ; 
   reg __394175_394175;
   reg _394176_394176 ; 
   reg __394176_394176;
   reg _394177_394177 ; 
   reg __394177_394177;
   reg _394178_394178 ; 
   reg __394178_394178;
   reg _394179_394179 ; 
   reg __394179_394179;
   reg _394180_394180 ; 
   reg __394180_394180;
   reg _394181_394181 ; 
   reg __394181_394181;
   reg _394182_394182 ; 
   reg __394182_394182;
   reg _394183_394183 ; 
   reg __394183_394183;
   reg _394184_394184 ; 
   reg __394184_394184;
   reg _394185_394185 ; 
   reg __394185_394185;
   reg _394186_394186 ; 
   reg __394186_394186;
   reg _394187_394187 ; 
   reg __394187_394187;
   reg _394188_394188 ; 
   reg __394188_394188;
   reg _394189_394189 ; 
   reg __394189_394189;
   reg _394190_394190 ; 
   reg __394190_394190;
   reg _394191_394191 ; 
   reg __394191_394191;
   reg _394192_394192 ; 
   reg __394192_394192;
   reg _394193_394193 ; 
   reg __394193_394193;
   reg _394194_394194 ; 
   reg __394194_394194;
   reg _394195_394195 ; 
   reg __394195_394195;
   reg _394196_394196 ; 
   reg __394196_394196;
   reg _394197_394197 ; 
   reg __394197_394197;
   reg _394198_394198 ; 
   reg __394198_394198;
   reg _394199_394199 ; 
   reg __394199_394199;
   reg _394200_394200 ; 
   reg __394200_394200;
   reg _394201_394201 ; 
   reg __394201_394201;
   reg _394202_394202 ; 
   reg __394202_394202;
   reg _394203_394203 ; 
   reg __394203_394203;
   reg _394204_394204 ; 
   reg __394204_394204;
   reg _394205_394205 ; 
   reg __394205_394205;
   reg _394206_394206 ; 
   reg __394206_394206;
   reg _394207_394207 ; 
   reg __394207_394207;
   reg _394208_394208 ; 
   reg __394208_394208;
   reg _394209_394209 ; 
   reg __394209_394209;
   reg _394210_394210 ; 
   reg __394210_394210;
   reg _394211_394211 ; 
   reg __394211_394211;
   reg _394212_394212 ; 
   reg __394212_394212;
   reg _394213_394213 ; 
   reg __394213_394213;
   reg _394214_394214 ; 
   reg __394214_394214;
   reg _394215_394215 ; 
   reg __394215_394215;
   reg _394216_394216 ; 
   reg __394216_394216;
   reg _394217_394217 ; 
   reg __394217_394217;
   reg _394218_394218 ; 
   reg __394218_394218;
   reg _394219_394219 ; 
   reg __394219_394219;
   reg _394220_394220 ; 
   reg __394220_394220;
   reg _394221_394221 ; 
   reg __394221_394221;
   reg _394222_394222 ; 
   reg __394222_394222;
   reg _394223_394223 ; 
   reg __394223_394223;
   reg _394224_394224 ; 
   reg __394224_394224;
   reg _394225_394225 ; 
   reg __394225_394225;
   reg _394226_394226 ; 
   reg __394226_394226;
   reg _394227_394227 ; 
   reg __394227_394227;
   reg _394228_394228 ; 
   reg __394228_394228;
   reg _394229_394229 ; 
   reg __394229_394229;
   reg _394230_394230 ; 
   reg __394230_394230;
   reg _394231_394231 ; 
   reg __394231_394231;
   reg _394232_394232 ; 
   reg __394232_394232;
   reg _394233_394233 ; 
   reg __394233_394233;
   reg _394234_394234 ; 
   reg __394234_394234;
   reg _394235_394235 ; 
   reg __394235_394235;
   reg _394236_394236 ; 
   reg __394236_394236;
   reg _394237_394237 ; 
   reg __394237_394237;
   reg _394238_394238 ; 
   reg __394238_394238;
   reg _394239_394239 ; 
   reg __394239_394239;
   reg _394240_394240 ; 
   reg __394240_394240;
   reg _394241_394241 ; 
   reg __394241_394241;
   reg _394242_394242 ; 
   reg __394242_394242;
   reg _394243_394243 ; 
   reg __394243_394243;
   reg _394244_394244 ; 
   reg __394244_394244;
   reg _394245_394245 ; 
   reg __394245_394245;
   reg _394246_394246 ; 
   reg __394246_394246;
   reg _394247_394247 ; 
   reg __394247_394247;
   reg _394248_394248 ; 
   reg __394248_394248;
   reg _394249_394249 ; 
   reg __394249_394249;
   reg _394250_394250 ; 
   reg __394250_394250;
   reg _394251_394251 ; 
   reg __394251_394251;
   reg _394252_394252 ; 
   reg __394252_394252;
   reg _394253_394253 ; 
   reg __394253_394253;
   reg _394254_394254 ; 
   reg __394254_394254;
   reg _394255_394255 ; 
   reg __394255_394255;
   reg _394256_394256 ; 
   reg __394256_394256;
   reg _394257_394257 ; 
   reg __394257_394257;
   reg _394258_394258 ; 
   reg __394258_394258;
   reg _394259_394259 ; 
   reg __394259_394259;
   reg _394260_394260 ; 
   reg __394260_394260;
   reg _394261_394261 ; 
   reg __394261_394261;
   reg _394262_394262 ; 
   reg __394262_394262;
   reg _394263_394263 ; 
   reg __394263_394263;
   reg _394264_394264 ; 
   reg __394264_394264;
   reg _394265_394265 ; 
   reg __394265_394265;
   reg _394266_394266 ; 
   reg __394266_394266;
   reg _394267_394267 ; 
   reg __394267_394267;
   reg _394268_394268 ; 
   reg __394268_394268;
   reg _394269_394269 ; 
   reg __394269_394269;
   reg _394270_394270 ; 
   reg __394270_394270;
   reg _394271_394271 ; 
   reg __394271_394271;
   reg _394272_394272 ; 
   reg __394272_394272;
   reg _394273_394273 ; 
   reg __394273_394273;
   reg _394274_394274 ; 
   reg __394274_394274;
   reg _394275_394275 ; 
   reg __394275_394275;
   reg _394276_394276 ; 
   reg __394276_394276;
   reg _394277_394277 ; 
   reg __394277_394277;
   reg _394278_394278 ; 
   reg __394278_394278;
   reg _394279_394279 ; 
   reg __394279_394279;
   reg _394280_394280 ; 
   reg __394280_394280;
   reg _394281_394281 ; 
   reg __394281_394281;
   reg _394282_394282 ; 
   reg __394282_394282;
   reg _394283_394283 ; 
   reg __394283_394283;
   reg _394284_394284 ; 
   reg __394284_394284;
   reg _394285_394285 ; 
   reg __394285_394285;
   reg _394286_394286 ; 
   reg __394286_394286;
   reg _394287_394287 ; 
   reg __394287_394287;
   reg _394288_394288 ; 
   reg __394288_394288;
   reg _394289_394289 ; 
   reg __394289_394289;
   reg _394290_394290 ; 
   reg __394290_394290;
   reg _394291_394291 ; 
   reg __394291_394291;
   reg _394292_394292 ; 
   reg __394292_394292;
   reg _394293_394293 ; 
   reg __394293_394293;
   reg _394294_394294 ; 
   reg __394294_394294;
   reg _394295_394295 ; 
   reg __394295_394295;
   reg _394296_394296 ; 
   reg __394296_394296;
   reg _394297_394297 ; 
   reg __394297_394297;
   reg _394298_394298 ; 
   reg __394298_394298;
   reg _394299_394299 ; 
   reg __394299_394299;
   reg _394300_394300 ; 
   reg __394300_394300;
   reg _394301_394301 ; 
   reg __394301_394301;
   reg _394302_394302 ; 
   reg __394302_394302;
   reg _394303_394303 ; 
   reg __394303_394303;
   reg _394304_394304 ; 
   reg __394304_394304;
   reg _394305_394305 ; 
   reg __394305_394305;
   reg _394306_394306 ; 
   reg __394306_394306;
   reg _394307_394307 ; 
   reg __394307_394307;
   reg _394308_394308 ; 
   reg __394308_394308;
   reg _394309_394309 ; 
   reg __394309_394309;
   reg _394310_394310 ; 
   reg __394310_394310;
   reg _394311_394311 ; 
   reg __394311_394311;
   reg _394312_394312 ; 
   reg __394312_394312;
   reg _394313_394313 ; 
   reg __394313_394313;
   reg _394314_394314 ; 
   reg __394314_394314;
   reg _394315_394315 ; 
   reg __394315_394315;
   reg _394316_394316 ; 
   reg __394316_394316;
   reg _394317_394317 ; 
   reg __394317_394317;
   reg _394318_394318 ; 
   reg __394318_394318;
   reg _394319_394319 ; 
   reg __394319_394319;
   reg _394320_394320 ; 
   reg __394320_394320;
   reg _394321_394321 ; 
   reg __394321_394321;
   reg _394322_394322 ; 
   reg __394322_394322;
   reg _394323_394323 ; 
   reg __394323_394323;
   reg _394324_394324 ; 
   reg __394324_394324;
   reg _394325_394325 ; 
   reg __394325_394325;
   reg _394326_394326 ; 
   reg __394326_394326;
   reg _394327_394327 ; 
   reg __394327_394327;
   reg _394328_394328 ; 
   reg __394328_394328;
   reg _394329_394329 ; 
   reg __394329_394329;
   reg _394330_394330 ; 
   reg __394330_394330;
   reg _394331_394331 ; 
   reg __394331_394331;
   reg _394332_394332 ; 
   reg __394332_394332;
   reg _394333_394333 ; 
   reg __394333_394333;
   reg _394334_394334 ; 
   reg __394334_394334;
   reg _394335_394335 ; 
   reg __394335_394335;
   reg _394336_394336 ; 
   reg __394336_394336;
   reg _394337_394337 ; 
   reg __394337_394337;
   reg _394338_394338 ; 
   reg __394338_394338;
   reg _394339_394339 ; 
   reg __394339_394339;
   reg _394340_394340 ; 
   reg __394340_394340;
   reg _394341_394341 ; 
   reg __394341_394341;
   reg _394342_394342 ; 
   reg __394342_394342;
   reg _394343_394343 ; 
   reg __394343_394343;
   reg _394344_394344 ; 
   reg __394344_394344;
   reg _394345_394345 ; 
   reg __394345_394345;
   reg _394346_394346 ; 
   reg __394346_394346;
   reg _394347_394347 ; 
   reg __394347_394347;
   reg _394348_394348 ; 
   reg __394348_394348;
   reg _394349_394349 ; 
   reg __394349_394349;
   reg _394350_394350 ; 
   reg __394350_394350;
   reg _394351_394351 ; 
   reg __394351_394351;
   reg _394352_394352 ; 
   reg __394352_394352;
   reg _394353_394353 ; 
   reg __394353_394353;
   reg _394354_394354 ; 
   reg __394354_394354;
   reg _394355_394355 ; 
   reg __394355_394355;
   reg _394356_394356 ; 
   reg __394356_394356;
   reg _394357_394357 ; 
   reg __394357_394357;
   reg _394358_394358 ; 
   reg __394358_394358;
   reg _394359_394359 ; 
   reg __394359_394359;
   reg _394360_394360 ; 
   reg __394360_394360;
   reg _394361_394361 ; 
   reg __394361_394361;
   reg _394362_394362 ; 
   reg __394362_394362;
   reg _394363_394363 ; 
   reg __394363_394363;
   reg _394364_394364 ; 
   reg __394364_394364;
   reg _394365_394365 ; 
   reg __394365_394365;
   reg _394366_394366 ; 
   reg __394366_394366;
   reg _394367_394367 ; 
   reg __394367_394367;
   reg _394368_394368 ; 
   reg __394368_394368;
   reg _394369_394369 ; 
   reg __394369_394369;
   reg _394370_394370 ; 
   reg __394370_394370;
   reg _394371_394371 ; 
   reg __394371_394371;
   reg _394372_394372 ; 
   reg __394372_394372;
   reg _394373_394373 ; 
   reg __394373_394373;
   reg _394374_394374 ; 
   reg __394374_394374;
   reg _394375_394375 ; 
   reg __394375_394375;
   reg _394376_394376 ; 
   reg __394376_394376;
   reg _394377_394377 ; 
   reg __394377_394377;
   reg _394378_394378 ; 
   reg __394378_394378;
   reg _394379_394379 ; 
   reg __394379_394379;
   reg _394380_394380 ; 
   reg __394380_394380;
   reg _394381_394381 ; 
   reg __394381_394381;
   reg _394382_394382 ; 
   reg __394382_394382;
   reg _394383_394383 ; 
   reg __394383_394383;
   reg _394384_394384 ; 
   reg __394384_394384;
   reg _394385_394385 ; 
   reg __394385_394385;
   reg _394386_394386 ; 
   reg __394386_394386;
   reg _394387_394387 ; 
   reg __394387_394387;
   reg _394388_394388 ; 
   reg __394388_394388;
   reg _394389_394389 ; 
   reg __394389_394389;
   reg _394390_394390 ; 
   reg __394390_394390;
   reg _394391_394391 ; 
   reg __394391_394391;
   reg _394392_394392 ; 
   reg __394392_394392;
   reg _394393_394393 ; 
   reg __394393_394393;
   reg _394394_394394 ; 
   reg __394394_394394;
   reg _394395_394395 ; 
   reg __394395_394395;
   reg _394396_394396 ; 
   reg __394396_394396;
   reg _394397_394397 ; 
   reg __394397_394397;
   reg _394398_394398 ; 
   reg __394398_394398;
   reg _394399_394399 ; 
   reg __394399_394399;
   reg _394400_394400 ; 
   reg __394400_394400;
   reg _394401_394401 ; 
   reg __394401_394401;
   reg _394402_394402 ; 
   reg __394402_394402;
   reg _394403_394403 ; 
   reg __394403_394403;
   reg _394404_394404 ; 
   reg __394404_394404;
   reg _394405_394405 ; 
   reg __394405_394405;
   reg _394406_394406 ; 
   reg __394406_394406;
   reg _394407_394407 ; 
   reg __394407_394407;
   reg _394408_394408 ; 
   reg __394408_394408;
   reg _394409_394409 ; 
   reg __394409_394409;
   reg _394410_394410 ; 
   reg __394410_394410;
   reg _394411_394411 ; 
   reg __394411_394411;
   reg _394412_394412 ; 
   reg __394412_394412;
   reg _394413_394413 ; 
   reg __394413_394413;
   reg _394414_394414 ; 
   reg __394414_394414;
   reg _394415_394415 ; 
   reg __394415_394415;
   reg _394416_394416 ; 
   reg __394416_394416;
   reg _394417_394417 ; 
   reg __394417_394417;
   reg _394418_394418 ; 
   reg __394418_394418;
   reg _394419_394419 ; 
   reg __394419_394419;
   reg _394420_394420 ; 
   reg __394420_394420;
   reg _394421_394421 ; 
   reg __394421_394421;
   reg _394422_394422 ; 
   reg __394422_394422;
   reg _394423_394423 ; 
   reg __394423_394423;
   reg _394424_394424 ; 
   reg __394424_394424;
   reg _394425_394425 ; 
   reg __394425_394425;
   reg _394426_394426 ; 
   reg __394426_394426;
   reg _394427_394427 ; 
   reg __394427_394427;
   reg _394428_394428 ; 
   reg __394428_394428;
   reg _394429_394429 ; 
   reg __394429_394429;
   reg _394430_394430 ; 
   reg __394430_394430;
   reg _394431_394431 ; 
   reg __394431_394431;
   reg _394432_394432 ; 
   reg __394432_394432;
   reg _394433_394433 ; 
   reg __394433_394433;
   reg _394434_394434 ; 
   reg __394434_394434;
   reg _394435_394435 ; 
   reg __394435_394435;
   reg _394436_394436 ; 
   reg __394436_394436;
   reg _394437_394437 ; 
   reg __394437_394437;
   reg _394438_394438 ; 
   reg __394438_394438;
   reg _394439_394439 ; 
   reg __394439_394439;
   reg _394440_394440 ; 
   reg __394440_394440;
   reg _394441_394441 ; 
   reg __394441_394441;
   reg _394442_394442 ; 
   reg __394442_394442;
   reg _394443_394443 ; 
   reg __394443_394443;
   reg _394444_394444 ; 
   reg __394444_394444;
   reg _394445_394445 ; 
   reg __394445_394445;
   reg _394446_394446 ; 
   reg __394446_394446;
   reg _394447_394447 ; 
   reg __394447_394447;
   reg _394448_394448 ; 
   reg __394448_394448;
   reg _394449_394449 ; 
   reg __394449_394449;
   reg _394450_394450 ; 
   reg __394450_394450;
   reg _394451_394451 ; 
   reg __394451_394451;
   reg _394452_394452 ; 
   reg __394452_394452;
   reg _394453_394453 ; 
   reg __394453_394453;
   reg _394454_394454 ; 
   reg __394454_394454;
   reg _394455_394455 ; 
   reg __394455_394455;
   reg _394456_394456 ; 
   reg __394456_394456;
   reg _394457_394457 ; 
   reg __394457_394457;
   reg _394458_394458 ; 
   reg __394458_394458;
   reg _394459_394459 ; 
   reg __394459_394459;
   reg _394460_394460 ; 
   reg __394460_394460;
   reg _394461_394461 ; 
   reg __394461_394461;
   reg _394462_394462 ; 
   reg __394462_394462;
   reg _394463_394463 ; 
   reg __394463_394463;
   reg _394464_394464 ; 
   reg __394464_394464;
   reg _394465_394465 ; 
   reg __394465_394465;
   reg _394466_394466 ; 
   reg __394466_394466;
   reg _394467_394467 ; 
   reg __394467_394467;
   reg _394468_394468 ; 
   reg __394468_394468;
   reg _394469_394469 ; 
   reg __394469_394469;
   reg _394470_394470 ; 
   reg __394470_394470;
   reg _394471_394471 ; 
   reg __394471_394471;
   reg _394472_394472 ; 
   reg __394472_394472;
   reg _394473_394473 ; 
   reg __394473_394473;
   reg _394474_394474 ; 
   reg __394474_394474;
   reg _394475_394475 ; 
   reg __394475_394475;
   reg _394476_394476 ; 
   reg __394476_394476;
   reg _394477_394477 ; 
   reg __394477_394477;
   reg _394478_394478 ; 
   reg __394478_394478;
   reg _394479_394479 ; 
   reg __394479_394479;
   reg _394480_394480 ; 
   reg __394480_394480;
   reg _394481_394481 ; 
   reg __394481_394481;
   reg _394482_394482 ; 
   reg __394482_394482;
   reg _394483_394483 ; 
   reg __394483_394483;
   reg _394484_394484 ; 
   reg __394484_394484;
   reg _394485_394485 ; 
   reg __394485_394485;
   reg _394486_394486 ; 
   reg __394486_394486;
   reg _394487_394487 ; 
   reg __394487_394487;
   reg _394488_394488 ; 
   reg __394488_394488;
   reg _394489_394489 ; 
   reg __394489_394489;
   reg _394490_394490 ; 
   reg __394490_394490;
   reg _394491_394491 ; 
   reg __394491_394491;
   reg _394492_394492 ; 
   reg __394492_394492;
   reg _394493_394493 ; 
   reg __394493_394493;
   reg _394494_394494 ; 
   reg __394494_394494;
   reg _394495_394495 ; 
   reg __394495_394495;
   reg _394496_394496 ; 
   reg __394496_394496;
   reg _394497_394497 ; 
   reg __394497_394497;
   reg _394498_394498 ; 
   reg __394498_394498;
   reg _394499_394499 ; 
   reg __394499_394499;
   reg _394500_394500 ; 
   reg __394500_394500;
   reg _394501_394501 ; 
   reg __394501_394501;
   reg _394502_394502 ; 
   reg __394502_394502;
   reg _394503_394503 ; 
   reg __394503_394503;
   reg _394504_394504 ; 
   reg __394504_394504;
   reg _394505_394505 ; 
   reg __394505_394505;
   reg _394506_394506 ; 
   reg __394506_394506;
   reg _394507_394507 ; 
   reg __394507_394507;
   reg _394508_394508 ; 
   reg __394508_394508;
   reg _394509_394509 ; 
   reg __394509_394509;
   reg _394510_394510 ; 
   reg __394510_394510;
   reg _394511_394511 ; 
   reg __394511_394511;
   reg _394512_394512 ; 
   reg __394512_394512;
   reg _394513_394513 ; 
   reg __394513_394513;
   reg _394514_394514 ; 
   reg __394514_394514;
   reg _394515_394515 ; 
   reg __394515_394515;
   reg _394516_394516 ; 
   reg __394516_394516;
   reg _394517_394517 ; 
   reg __394517_394517;
   reg _394518_394518 ; 
   reg __394518_394518;
   reg _394519_394519 ; 
   reg __394519_394519;
   reg _394520_394520 ; 
   reg __394520_394520;
   reg _394521_394521 ; 
   reg __394521_394521;
   reg _394522_394522 ; 
   reg __394522_394522;
   reg _394523_394523 ; 
   reg __394523_394523;
   reg _394524_394524 ; 
   reg __394524_394524;
   reg _394525_394525 ; 
   reg __394525_394525;
   reg _394526_394526 ; 
   reg __394526_394526;
   reg _394527_394527 ; 
   reg __394527_394527;
   reg _394528_394528 ; 
   reg __394528_394528;
   reg _394529_394529 ; 
   reg __394529_394529;
   reg _394530_394530 ; 
   reg __394530_394530;
   reg _394531_394531 ; 
   reg __394531_394531;
   reg _394532_394532 ; 
   reg __394532_394532;
   reg _394533_394533 ; 
   reg __394533_394533;
   reg _394534_394534 ; 
   reg __394534_394534;
   reg _394535_394535 ; 
   reg __394535_394535;
   reg _394536_394536 ; 
   reg __394536_394536;
   reg _394537_394537 ; 
   reg __394537_394537;
   reg _394538_394538 ; 
   reg __394538_394538;
   reg _394539_394539 ; 
   reg __394539_394539;
   reg _394540_394540 ; 
   reg __394540_394540;
   reg _394541_394541 ; 
   reg __394541_394541;
   reg _394542_394542 ; 
   reg __394542_394542;
   reg _394543_394543 ; 
   reg __394543_394543;
   reg _394544_394544 ; 
   reg __394544_394544;
   reg _394545_394545 ; 
   reg __394545_394545;
   reg _394546_394546 ; 
   reg __394546_394546;
   reg _394547_394547 ; 
   reg __394547_394547;
   reg _394548_394548 ; 
   reg __394548_394548;
   reg _394549_394549 ; 
   reg __394549_394549;
   reg _394550_394550 ; 
   reg __394550_394550;
   reg _394551_394551 ; 
   reg __394551_394551;
   reg _394552_394552 ; 
   reg __394552_394552;
   reg _394553_394553 ; 
   reg __394553_394553;
   reg _394554_394554 ; 
   reg __394554_394554;
   reg _394555_394555 ; 
   reg __394555_394555;
   reg _394556_394556 ; 
   reg __394556_394556;
   reg _394557_394557 ; 
   reg __394557_394557;
   reg _394558_394558 ; 
   reg __394558_394558;
   reg _394559_394559 ; 
   reg __394559_394559;
   reg _394560_394560 ; 
   reg __394560_394560;
   reg _394561_394561 ; 
   reg __394561_394561;
   reg _394562_394562 ; 
   reg __394562_394562;
   reg _394563_394563 ; 
   reg __394563_394563;
   reg _394564_394564 ; 
   reg __394564_394564;
   reg _394565_394565 ; 
   reg __394565_394565;
   reg _394566_394566 ; 
   reg __394566_394566;
   reg _394567_394567 ; 
   reg __394567_394567;
   reg _394568_394568 ; 
   reg __394568_394568;
   reg _394569_394569 ; 
   reg __394569_394569;
   reg _394570_394570 ; 
   reg __394570_394570;
   reg _394571_394571 ; 
   reg __394571_394571;
   reg _394572_394572 ; 
   reg __394572_394572;
   reg _394573_394573 ; 
   reg __394573_394573;
   reg _394574_394574 ; 
   reg __394574_394574;
   reg _394575_394575 ; 
   reg __394575_394575;
   reg _394576_394576 ; 
   reg __394576_394576;
   reg _394577_394577 ; 
   reg __394577_394577;
   reg _394578_394578 ; 
   reg __394578_394578;
   reg _394579_394579 ; 
   reg __394579_394579;
   reg _394580_394580 ; 
   reg __394580_394580;
   reg _394581_394581 ; 
   reg __394581_394581;
   reg _394582_394582 ; 
   reg __394582_394582;
   reg _394583_394583 ; 
   reg __394583_394583;
   reg _394584_394584 ; 
   reg __394584_394584;
   reg _394585_394585 ; 
   reg __394585_394585;
   reg _394586_394586 ; 
   reg __394586_394586;
   reg _394587_394587 ; 
   reg __394587_394587;
   reg _394588_394588 ; 
   reg __394588_394588;
   reg _394589_394589 ; 
   reg __394589_394589;
   reg _394590_394590 ; 
   reg __394590_394590;
   reg _394591_394591 ; 
   reg __394591_394591;
   reg _394592_394592 ; 
   reg __394592_394592;
   reg _394593_394593 ; 
   reg __394593_394593;
   reg _394594_394594 ; 
   reg __394594_394594;
   reg _394595_394595 ; 
   reg __394595_394595;
   reg _394596_394596 ; 
   reg __394596_394596;
   reg _394597_394597 ; 
   reg __394597_394597;
   reg _394598_394598 ; 
   reg __394598_394598;
   reg _394599_394599 ; 
   reg __394599_394599;
   reg _394600_394600 ; 
   reg __394600_394600;
   reg _394601_394601 ; 
   reg __394601_394601;
   reg _394602_394602 ; 
   reg __394602_394602;
   reg _394603_394603 ; 
   reg __394603_394603;
   reg _394604_394604 ; 
   reg __394604_394604;
   reg _394605_394605 ; 
   reg __394605_394605;
   reg _394606_394606 ; 
   reg __394606_394606;
   reg _394607_394607 ; 
   reg __394607_394607;
   reg _394608_394608 ; 
   reg __394608_394608;
   reg _394609_394609 ; 
   reg __394609_394609;
   reg _394610_394610 ; 
   reg __394610_394610;
   reg _394611_394611 ; 
   reg __394611_394611;
   reg _394612_394612 ; 
   reg __394612_394612;
   reg _394613_394613 ; 
   reg __394613_394613;
   reg _394614_394614 ; 
   reg __394614_394614;
   reg _394615_394615 ; 
   reg __394615_394615;
   reg _394616_394616 ; 
   reg __394616_394616;
   reg _394617_394617 ; 
   reg __394617_394617;
   reg _394618_394618 ; 
   reg __394618_394618;
   reg _394619_394619 ; 
   reg __394619_394619;
   reg _394620_394620 ; 
   reg __394620_394620;
   reg _394621_394621 ; 
   reg __394621_394621;
   reg _394622_394622 ; 
   reg __394622_394622;
   reg _394623_394623 ; 
   reg __394623_394623;
   reg _394624_394624 ; 
   reg __394624_394624;
   reg _394625_394625 ; 
   reg __394625_394625;
   reg _394626_394626 ; 
   reg __394626_394626;
   reg _394627_394627 ; 
   reg __394627_394627;
   reg _394628_394628 ; 
   reg __394628_394628;
   reg _394629_394629 ; 
   reg __394629_394629;
   reg _394630_394630 ; 
   reg __394630_394630;
   reg _394631_394631 ; 
   reg __394631_394631;
   reg _394632_394632 ; 
   reg __394632_394632;
   reg _394633_394633 ; 
   reg __394633_394633;
   reg _394634_394634 ; 
   reg __394634_394634;
   reg _394635_394635 ; 
   reg __394635_394635;
   reg _394636_394636 ; 
   reg __394636_394636;
   reg _394637_394637 ; 
   reg __394637_394637;
   reg _394638_394638 ; 
   reg __394638_394638;
   reg _394639_394639 ; 
   reg __394639_394639;
   reg _394640_394640 ; 
   reg __394640_394640;
   reg _394641_394641 ; 
   reg __394641_394641;
   reg _394642_394642 ; 
   reg __394642_394642;
   reg _394643_394643 ; 
   reg __394643_394643;
   reg _394644_394644 ; 
   reg __394644_394644;
   reg _394645_394645 ; 
   reg __394645_394645;
   reg _394646_394646 ; 
   reg __394646_394646;
   reg _394647_394647 ; 
   reg __394647_394647;
   reg _394648_394648 ; 
   reg __394648_394648;
   reg _394649_394649 ; 
   reg __394649_394649;
   reg _394650_394650 ; 
   reg __394650_394650;
   reg _394651_394651 ; 
   reg __394651_394651;
   reg _394652_394652 ; 
   reg __394652_394652;
   reg _394653_394653 ; 
   reg __394653_394653;
   reg _394654_394654 ; 
   reg __394654_394654;
   reg _394655_394655 ; 
   reg __394655_394655;
   reg _394656_394656 ; 
   reg __394656_394656;
   reg _394657_394657 ; 
   reg __394657_394657;
   reg _394658_394658 ; 
   reg __394658_394658;
   reg _394659_394659 ; 
   reg __394659_394659;
   reg _394660_394660 ; 
   reg __394660_394660;
   reg _394661_394661 ; 
   reg __394661_394661;
   reg _394662_394662 ; 
   reg __394662_394662;
   reg _394663_394663 ; 
   reg __394663_394663;
   reg _394664_394664 ; 
   reg __394664_394664;
   reg _394665_394665 ; 
   reg __394665_394665;
   reg _394666_394666 ; 
   reg __394666_394666;
   reg _394667_394667 ; 
   reg __394667_394667;
   reg _394668_394668 ; 
   reg __394668_394668;
   reg _394669_394669 ; 
   reg __394669_394669;
   reg _394670_394670 ; 
   reg __394670_394670;
   reg _394671_394671 ; 
   reg __394671_394671;
   reg _394672_394672 ; 
   reg __394672_394672;
   reg _394673_394673 ; 
   reg __394673_394673;
   reg _394674_394674 ; 
   reg __394674_394674;
   reg _394675_394675 ; 
   reg __394675_394675;
   reg _394676_394676 ; 
   reg __394676_394676;
   reg _394677_394677 ; 
   reg __394677_394677;
   reg _394678_394678 ; 
   reg __394678_394678;
   reg _394679_394679 ; 
   reg __394679_394679;
   reg _394680_394680 ; 
   reg __394680_394680;
   reg _394681_394681 ; 
   reg __394681_394681;
   reg _394682_394682 ; 
   reg __394682_394682;
   reg _394683_394683 ; 
   reg __394683_394683;
   reg _394684_394684 ; 
   reg __394684_394684;
   reg _394685_394685 ; 
   reg __394685_394685;
   reg _394686_394686 ; 
   reg __394686_394686;
   reg _394687_394687 ; 
   reg __394687_394687;
   reg _394688_394688 ; 
   reg __394688_394688;
   reg _394689_394689 ; 
   reg __394689_394689;
   reg _394690_394690 ; 
   reg __394690_394690;
   reg _394691_394691 ; 
   reg __394691_394691;
   reg _394692_394692 ; 
   reg __394692_394692;
   reg _394693_394693 ; 
   reg __394693_394693;
   reg _394694_394694 ; 
   reg __394694_394694;
   reg _394695_394695 ; 
   reg __394695_394695;
   reg _394696_394696 ; 
   reg __394696_394696;
   reg _394697_394697 ; 
   reg __394697_394697;
   reg _394698_394698 ; 
   reg __394698_394698;
   reg _394699_394699 ; 
   reg __394699_394699;
   reg _394700_394700 ; 
   reg __394700_394700;
   reg _394701_394701 ; 
   reg __394701_394701;
   reg _394702_394702 ; 
   reg __394702_394702;
   reg _394703_394703 ; 
   reg __394703_394703;
   reg _394704_394704 ; 
   reg __394704_394704;
   reg _394705_394705 ; 
   reg __394705_394705;
   reg _394706_394706 ; 
   reg __394706_394706;
   reg _394707_394707 ; 
   reg __394707_394707;
   reg _394708_394708 ; 
   reg __394708_394708;
   reg _394709_394709 ; 
   reg __394709_394709;
   reg _394710_394710 ; 
   reg __394710_394710;
   reg _394711_394711 ; 
   reg __394711_394711;
   reg _394712_394712 ; 
   reg __394712_394712;
   reg _394713_394713 ; 
   reg __394713_394713;
   reg _394714_394714 ; 
   reg __394714_394714;
   reg _394715_394715 ; 
   reg __394715_394715;
   reg _394716_394716 ; 
   reg __394716_394716;
   reg _394717_394717 ; 
   reg __394717_394717;
   reg _394718_394718 ; 
   reg __394718_394718;
   reg _394719_394719 ; 
   reg __394719_394719;
   reg _394720_394720 ; 
   reg __394720_394720;
   reg _394721_394721 ; 
   reg __394721_394721;
   reg _394722_394722 ; 
   reg __394722_394722;
   reg _394723_394723 ; 
   reg __394723_394723;
   reg _394724_394724 ; 
   reg __394724_394724;
   reg _394725_394725 ; 
   reg __394725_394725;
   reg _394726_394726 ; 
   reg __394726_394726;
   reg _394727_394727 ; 
   reg __394727_394727;
   reg _394728_394728 ; 
   reg __394728_394728;
   reg _394729_394729 ; 
   reg __394729_394729;
   reg _394730_394730 ; 
   reg __394730_394730;
   reg _394731_394731 ; 
   reg __394731_394731;
   reg _394732_394732 ; 
   reg __394732_394732;
   reg _394733_394733 ; 
   reg __394733_394733;
   reg _394734_394734 ; 
   reg __394734_394734;
   reg _394735_394735 ; 
   reg __394735_394735;
   reg _394736_394736 ; 
   reg __394736_394736;
   reg _394737_394737 ; 
   reg __394737_394737;
   reg _394738_394738 ; 
   reg __394738_394738;
   reg _394739_394739 ; 
   reg __394739_394739;
   reg _394740_394740 ; 
   reg __394740_394740;
   reg _394741_394741 ; 
   reg __394741_394741;
   reg _394742_394742 ; 
   reg __394742_394742;
   reg _394743_394743 ; 
   reg __394743_394743;
   reg _394744_394744 ; 
   reg __394744_394744;
   reg _394745_394745 ; 
   reg __394745_394745;
   reg _394746_394746 ; 
   reg __394746_394746;
   reg _394747_394747 ; 
   reg __394747_394747;
   reg _394748_394748 ; 
   reg __394748_394748;
   reg _394749_394749 ; 
   reg __394749_394749;
   reg _394750_394750 ; 
   reg __394750_394750;
   reg _394751_394751 ; 
   reg __394751_394751;
   reg _394752_394752 ; 
   reg __394752_394752;
   reg _394753_394753 ; 
   reg __394753_394753;
   reg _394754_394754 ; 
   reg __394754_394754;
   reg _394755_394755 ; 
   reg __394755_394755;
   reg _394756_394756 ; 
   reg __394756_394756;
   reg _394757_394757 ; 
   reg __394757_394757;
   reg _394758_394758 ; 
   reg __394758_394758;
   reg _394759_394759 ; 
   reg __394759_394759;
   reg _394760_394760 ; 
   reg __394760_394760;
   reg _394761_394761 ; 
   reg __394761_394761;
   reg _394762_394762 ; 
   reg __394762_394762;
   reg _394763_394763 ; 
   reg __394763_394763;
   reg _394764_394764 ; 
   reg __394764_394764;
   reg _394765_394765 ; 
   reg __394765_394765;
   reg _394766_394766 ; 
   reg __394766_394766;
   reg _394767_394767 ; 
   reg __394767_394767;
   reg _394768_394768 ; 
   reg __394768_394768;
   reg _394769_394769 ; 
   reg __394769_394769;
   reg _394770_394770 ; 
   reg __394770_394770;
   reg _394771_394771 ; 
   reg __394771_394771;
   reg _394772_394772 ; 
   reg __394772_394772;
   reg _394773_394773 ; 
   reg __394773_394773;
   reg _394774_394774 ; 
   reg __394774_394774;
   reg _394775_394775 ; 
   reg __394775_394775;
   reg _394776_394776 ; 
   reg __394776_394776;
   reg _394777_394777 ; 
   reg __394777_394777;
   reg _394778_394778 ; 
   reg __394778_394778;
   reg _394779_394779 ; 
   reg __394779_394779;
   reg _394780_394780 ; 
   reg __394780_394780;
   reg _394781_394781 ; 
   reg __394781_394781;
   reg _394782_394782 ; 
   reg __394782_394782;
   reg _394783_394783 ; 
   reg __394783_394783;
   reg _394784_394784 ; 
   reg __394784_394784;
   reg _394785_394785 ; 
   reg __394785_394785;
   reg _394786_394786 ; 
   reg __394786_394786;
   reg _394787_394787 ; 
   reg __394787_394787;
   reg _394788_394788 ; 
   reg __394788_394788;
   reg _394789_394789 ; 
   reg __394789_394789;
   reg _394790_394790 ; 
   reg __394790_394790;
   reg _394791_394791 ; 
   reg __394791_394791;
   reg _394792_394792 ; 
   reg __394792_394792;
   reg _394793_394793 ; 
   reg __394793_394793;
   reg _394794_394794 ; 
   reg __394794_394794;
   reg _394795_394795 ; 
   reg __394795_394795;
   reg _394796_394796 ; 
   reg __394796_394796;
   reg _394797_394797 ; 
   reg __394797_394797;
   reg _394798_394798 ; 
   reg __394798_394798;
   reg _394799_394799 ; 
   reg __394799_394799;
   reg _394800_394800 ; 
   reg __394800_394800;
   reg _394801_394801 ; 
   reg __394801_394801;
   reg _394802_394802 ; 
   reg __394802_394802;
   reg _394803_394803 ; 
   reg __394803_394803;
   reg _394804_394804 ; 
   reg __394804_394804;
   reg _394805_394805 ; 
   reg __394805_394805;
   reg _394806_394806 ; 
   reg __394806_394806;
   reg _394807_394807 ; 
   reg __394807_394807;
   reg _394808_394808 ; 
   reg __394808_394808;
   reg _394809_394809 ; 
   reg __394809_394809;
   reg _394810_394810 ; 
   reg __394810_394810;
   reg _394811_394811 ; 
   reg __394811_394811;
   reg _394812_394812 ; 
   reg __394812_394812;
   reg _394813_394813 ; 
   reg __394813_394813;
   reg _394814_394814 ; 
   reg __394814_394814;
   reg _394815_394815 ; 
   reg __394815_394815;
   reg _394816_394816 ; 
   reg __394816_394816;
   reg _394817_394817 ; 
   reg __394817_394817;
   reg _394818_394818 ; 
   reg __394818_394818;
   reg _394819_394819 ; 
   reg __394819_394819;
   reg _394820_394820 ; 
   reg __394820_394820;
   reg _394821_394821 ; 
   reg __394821_394821;
   reg _394822_394822 ; 
   reg __394822_394822;
   reg _394823_394823 ; 
   reg __394823_394823;
   reg _394824_394824 ; 
   reg __394824_394824;
   reg _394825_394825 ; 
   reg __394825_394825;
   reg _394826_394826 ; 
   reg __394826_394826;
   reg _394827_394827 ; 
   reg __394827_394827;
   reg _394828_394828 ; 
   reg __394828_394828;
   reg _394829_394829 ; 
   reg __394829_394829;
   reg _394830_394830 ; 
   reg __394830_394830;
   reg _394831_394831 ; 
   reg __394831_394831;
   reg _394832_394832 ; 
   reg __394832_394832;
   reg _394833_394833 ; 
   reg __394833_394833;
   reg _394834_394834 ; 
   reg __394834_394834;
   reg _394835_394835 ; 
   reg __394835_394835;
   reg _394836_394836 ; 
   reg __394836_394836;
   reg _394837_394837 ; 
   reg __394837_394837;
   reg _394838_394838 ; 
   reg __394838_394838;
   reg _394839_394839 ; 
   reg __394839_394839;
   reg _394840_394840 ; 
   reg __394840_394840;
   reg _394841_394841 ; 
   reg __394841_394841;
   reg _394842_394842 ; 
   reg __394842_394842;
   reg _394843_394843 ; 
   reg __394843_394843;
   reg _394844_394844 ; 
   reg __394844_394844;
   reg _394845_394845 ; 
   reg __394845_394845;
   reg _394846_394846 ; 
   reg __394846_394846;
   reg _394847_394847 ; 
   reg __394847_394847;
   reg _394848_394848 ; 
   reg __394848_394848;
   reg _394849_394849 ; 
   reg __394849_394849;
   reg _394850_394850 ; 
   reg __394850_394850;
   reg _394851_394851 ; 
   reg __394851_394851;
   reg _394852_394852 ; 
   reg __394852_394852;
   reg _394853_394853 ; 
   reg __394853_394853;
   reg _394854_394854 ; 
   reg __394854_394854;
   reg _394855_394855 ; 
   reg __394855_394855;
   reg _394856_394856 ; 
   reg __394856_394856;
   reg _394857_394857 ; 
   reg __394857_394857;
   reg _394858_394858 ; 
   reg __394858_394858;
   reg _394859_394859 ; 
   reg __394859_394859;
   reg _394860_394860 ; 
   reg __394860_394860;
   reg _394861_394861 ; 
   reg __394861_394861;
   reg _394862_394862 ; 
   reg __394862_394862;
   reg _394863_394863 ; 
   reg __394863_394863;
   reg _394864_394864 ; 
   reg __394864_394864;
   reg _394865_394865 ; 
   reg __394865_394865;
   reg _394866_394866 ; 
   reg __394866_394866;
   reg _394867_394867 ; 
   reg __394867_394867;
   reg _394868_394868 ; 
   reg __394868_394868;
   reg _394869_394869 ; 
   reg __394869_394869;
   reg _394870_394870 ; 
   reg __394870_394870;
   reg _394871_394871 ; 
   reg __394871_394871;
   reg _394872_394872 ; 
   reg __394872_394872;
   reg _394873_394873 ; 
   reg __394873_394873;
   reg _394874_394874 ; 
   reg __394874_394874;
   reg _394875_394875 ; 
   reg __394875_394875;
   reg _394876_394876 ; 
   reg __394876_394876;
   reg _394877_394877 ; 
   reg __394877_394877;
   reg _394878_394878 ; 
   reg __394878_394878;
   reg _394879_394879 ; 
   reg __394879_394879;
   reg _394880_394880 ; 
   reg __394880_394880;
   reg _394881_394881 ; 
   reg __394881_394881;
   reg _394882_394882 ; 
   reg __394882_394882;
   reg _394883_394883 ; 
   reg __394883_394883;
   reg _394884_394884 ; 
   reg __394884_394884;
   reg _394885_394885 ; 
   reg __394885_394885;
   reg _394886_394886 ; 
   reg __394886_394886;
   reg _394887_394887 ; 
   reg __394887_394887;
   reg _394888_394888 ; 
   reg __394888_394888;
   reg _394889_394889 ; 
   reg __394889_394889;
   reg _394890_394890 ; 
   reg __394890_394890;
   reg _394891_394891 ; 
   reg __394891_394891;
   reg _394892_394892 ; 
   reg __394892_394892;
   reg _394893_394893 ; 
   reg __394893_394893;
   reg _394894_394894 ; 
   reg __394894_394894;
   reg _394895_394895 ; 
   reg __394895_394895;
   reg _394896_394896 ; 
   reg __394896_394896;
   reg _394897_394897 ; 
   reg __394897_394897;
   reg _394898_394898 ; 
   reg __394898_394898;
   reg _394899_394899 ; 
   reg __394899_394899;
   reg _394900_394900 ; 
   reg __394900_394900;
   reg _394901_394901 ; 
   reg __394901_394901;
   reg _394902_394902 ; 
   reg __394902_394902;
   reg _394903_394903 ; 
   reg __394903_394903;
   reg _394904_394904 ; 
   reg __394904_394904;
   reg _394905_394905 ; 
   reg __394905_394905;
   reg _394906_394906 ; 
   reg __394906_394906;
   reg _394907_394907 ; 
   reg __394907_394907;
   reg _394908_394908 ; 
   reg __394908_394908;
   reg _394909_394909 ; 
   reg __394909_394909;
   reg _394910_394910 ; 
   reg __394910_394910;
   reg _394911_394911 ; 
   reg __394911_394911;
   reg _394912_394912 ; 
   reg __394912_394912;
   reg _394913_394913 ; 
   reg __394913_394913;
   reg _394914_394914 ; 
   reg __394914_394914;
   reg _394915_394915 ; 
   reg __394915_394915;
   reg _394916_394916 ; 
   reg __394916_394916;
   reg _394917_394917 ; 
   reg __394917_394917;
   reg _394918_394918 ; 
   reg __394918_394918;
   reg _394919_394919 ; 
   reg __394919_394919;
   reg _394920_394920 ; 
   reg __394920_394920;
   reg _394921_394921 ; 
   reg __394921_394921;
   reg _394922_394922 ; 
   reg __394922_394922;
   reg _394923_394923 ; 
   reg __394923_394923;
   reg _394924_394924 ; 
   reg __394924_394924;
   reg _394925_394925 ; 
   reg __394925_394925;
   reg _394926_394926 ; 
   reg __394926_394926;
   reg _394927_394927 ; 
   reg __394927_394927;
   reg _394928_394928 ; 
   reg __394928_394928;
   reg _394929_394929 ; 
   reg __394929_394929;
   reg _394930_394930 ; 
   reg __394930_394930;
   reg _394931_394931 ; 
   reg __394931_394931;
   reg _394932_394932 ; 
   reg __394932_394932;
   reg _394933_394933 ; 
   reg __394933_394933;
   reg _394934_394934 ; 
   reg __394934_394934;
   reg _394935_394935 ; 
   reg __394935_394935;
   reg _394936_394936 ; 
   reg __394936_394936;
   reg _394937_394937 ; 
   reg __394937_394937;
   reg _394938_394938 ; 
   reg __394938_394938;
   reg _394939_394939 ; 
   reg __394939_394939;
   reg _394940_394940 ; 
   reg __394940_394940;
   reg _394941_394941 ; 
   reg __394941_394941;
   reg _394942_394942 ; 
   reg __394942_394942;
   reg _394943_394943 ; 
   reg __394943_394943;
   reg _394944_394944 ; 
   reg __394944_394944;
   reg _394945_394945 ; 
   reg __394945_394945;
   reg _394946_394946 ; 
   reg __394946_394946;
   reg _394947_394947 ; 
   reg __394947_394947;
   reg _394948_394948 ; 
   reg __394948_394948;
   reg _394949_394949 ; 
   reg __394949_394949;
   reg _394950_394950 ; 
   reg __394950_394950;
   reg _394951_394951 ; 
   reg __394951_394951;
   reg _394952_394952 ; 
   reg __394952_394952;
   reg _394953_394953 ; 
   reg __394953_394953;
   reg _394954_394954 ; 
   reg __394954_394954;
   reg _394955_394955 ; 
   reg __394955_394955;
   reg _394956_394956 ; 
   reg __394956_394956;
   reg _394957_394957 ; 
   reg __394957_394957;
   reg _394958_394958 ; 
   reg __394958_394958;
   reg _394959_394959 ; 
   reg __394959_394959;
   reg _394960_394960 ; 
   reg __394960_394960;
   reg _394961_394961 ; 
   reg __394961_394961;
   reg _394962_394962 ; 
   reg __394962_394962;
   reg _394963_394963 ; 
   reg __394963_394963;
   reg _394964_394964 ; 
   reg __394964_394964;
   reg _394965_394965 ; 
   reg __394965_394965;
   reg _394966_394966 ; 
   reg __394966_394966;
   reg _394967_394967 ; 
   reg __394967_394967;
   reg _394968_394968 ; 
   reg __394968_394968;
   reg _394969_394969 ; 
   reg __394969_394969;
   reg _394970_394970 ; 
   reg __394970_394970;
   reg _394971_394971 ; 
   reg __394971_394971;
   reg _394972_394972 ; 
   reg __394972_394972;
   reg _394973_394973 ; 
   reg __394973_394973;
   reg _394974_394974 ; 
   reg __394974_394974;
   reg _394975_394975 ; 
   reg __394975_394975;
   reg _394976_394976 ; 
   reg __394976_394976;
   reg _394977_394977 ; 
   reg __394977_394977;
   reg _394978_394978 ; 
   reg __394978_394978;
   reg _394979_394979 ; 
   reg __394979_394979;
   reg _394980_394980 ; 
   reg __394980_394980;
   reg _394981_394981 ; 
   reg __394981_394981;
   reg _394982_394982 ; 
   reg __394982_394982;
   reg _394983_394983 ; 
   reg __394983_394983;
   reg _394984_394984 ; 
   reg __394984_394984;
   reg _394985_394985 ; 
   reg __394985_394985;
   reg _394986_394986 ; 
   reg __394986_394986;
   reg _394987_394987 ; 
   reg __394987_394987;
   reg _394988_394988 ; 
   reg __394988_394988;
   reg _394989_394989 ; 
   reg __394989_394989;
   reg _394990_394990 ; 
   reg __394990_394990;
   reg _394991_394991 ; 
   reg __394991_394991;
   reg _394992_394992 ; 
   reg __394992_394992;
   reg _394993_394993 ; 
   reg __394993_394993;
   reg _394994_394994 ; 
   reg __394994_394994;
   reg _394995_394995 ; 
   reg __394995_394995;
   reg _394996_394996 ; 
   reg __394996_394996;
   reg _394997_394997 ; 
   reg __394997_394997;
   reg _394998_394998 ; 
   reg __394998_394998;
   reg _394999_394999 ; 
   reg __394999_394999;
   reg _395000_395000 ; 
   reg __395000_395000;
   reg _395001_395001 ; 
   reg __395001_395001;
   reg _395002_395002 ; 
   reg __395002_395002;
   reg _395003_395003 ; 
   reg __395003_395003;
   reg _395004_395004 ; 
   reg __395004_395004;
   reg _395005_395005 ; 
   reg __395005_395005;
   reg _395006_395006 ; 
   reg __395006_395006;
   reg _395007_395007 ; 
   reg __395007_395007;
   reg _395008_395008 ; 
   reg __395008_395008;
   reg _395009_395009 ; 
   reg __395009_395009;
   reg _395010_395010 ; 
   reg __395010_395010;
   reg _395011_395011 ; 
   reg __395011_395011;
   reg _395012_395012 ; 
   reg __395012_395012;
   reg _395013_395013 ; 
   reg __395013_395013;
   reg _395014_395014 ; 
   reg __395014_395014;
   reg _395015_395015 ; 
   reg __395015_395015;
   reg _395016_395016 ; 
   reg __395016_395016;
   reg _395017_395017 ; 
   reg __395017_395017;
   reg _395018_395018 ; 
   reg __395018_395018;
   reg _395019_395019 ; 
   reg __395019_395019;
   reg _395020_395020 ; 
   reg __395020_395020;
   reg _395021_395021 ; 
   reg __395021_395021;
   reg _395022_395022 ; 
   reg __395022_395022;
   reg _395023_395023 ; 
   reg __395023_395023;
   reg _395024_395024 ; 
   reg __395024_395024;
   reg _395025_395025 ; 
   reg __395025_395025;
   reg _395026_395026 ; 
   reg __395026_395026;
   reg _395027_395027 ; 
   reg __395027_395027;
   reg _395028_395028 ; 
   reg __395028_395028;
   reg _395029_395029 ; 
   reg __395029_395029;
   reg _395030_395030 ; 
   reg __395030_395030;
   reg _395031_395031 ; 
   reg __395031_395031;
   reg _395032_395032 ; 
   reg __395032_395032;
   reg _395033_395033 ; 
   reg __395033_395033;
   reg _395034_395034 ; 
   reg __395034_395034;
   reg _395035_395035 ; 
   reg __395035_395035;
   reg _395036_395036 ; 
   reg __395036_395036;
   reg _395037_395037 ; 
   reg __395037_395037;
   reg _395038_395038 ; 
   reg __395038_395038;
   reg _395039_395039 ; 
   reg __395039_395039;
   reg _395040_395040 ; 
   reg __395040_395040;
   reg _395041_395041 ; 
   reg __395041_395041;
   reg _395042_395042 ; 
   reg __395042_395042;
   reg _395043_395043 ; 
   reg __395043_395043;
   reg _395044_395044 ; 
   reg __395044_395044;
   reg _395045_395045 ; 
   reg __395045_395045;
   reg _395046_395046 ; 
   reg __395046_395046;
   reg _395047_395047 ; 
   reg __395047_395047;
   reg _395048_395048 ; 
   reg __395048_395048;
   reg _395049_395049 ; 
   reg __395049_395049;
   reg _395050_395050 ; 
   reg __395050_395050;
   reg _395051_395051 ; 
   reg __395051_395051;
   reg _395052_395052 ; 
   reg __395052_395052;
   reg _395053_395053 ; 
   reg __395053_395053;
   reg _395054_395054 ; 
   reg __395054_395054;
   reg _395055_395055 ; 
   reg __395055_395055;
   reg _395056_395056 ; 
   reg __395056_395056;
   reg _395057_395057 ; 
   reg __395057_395057;
   reg _395058_395058 ; 
   reg __395058_395058;
   reg _395059_395059 ; 
   reg __395059_395059;
   reg _395060_395060 ; 
   reg __395060_395060;
   reg _395061_395061 ; 
   reg __395061_395061;
   reg _395062_395062 ; 
   reg __395062_395062;
   reg _395063_395063 ; 
   reg __395063_395063;
   reg _395064_395064 ; 
   reg __395064_395064;
   reg _395065_395065 ; 
   reg __395065_395065;
   reg _395066_395066 ; 
   reg __395066_395066;
   reg _395067_395067 ; 
   reg __395067_395067;
   reg _395068_395068 ; 
   reg __395068_395068;
   reg _395069_395069 ; 
   reg __395069_395069;
   reg _395070_395070 ; 
   reg __395070_395070;
   reg _395071_395071 ; 
   reg __395071_395071;
   reg _395072_395072 ; 
   reg __395072_395072;
   reg _395073_395073 ; 
   reg __395073_395073;
   reg _395074_395074 ; 
   reg __395074_395074;
   reg _395075_395075 ; 
   reg __395075_395075;
   reg _395076_395076 ; 
   reg __395076_395076;
   reg _395077_395077 ; 
   reg __395077_395077;
   reg _395078_395078 ; 
   reg __395078_395078;
   reg _395079_395079 ; 
   reg __395079_395079;
   reg _395080_395080 ; 
   reg __395080_395080;
   reg _395081_395081 ; 
   reg __395081_395081;
   reg _395082_395082 ; 
   reg __395082_395082;
   reg _395083_395083 ; 
   reg __395083_395083;
   reg _395084_395084 ; 
   reg __395084_395084;
   reg _395085_395085 ; 
   reg __395085_395085;
   reg _395086_395086 ; 
   reg __395086_395086;
   reg _395087_395087 ; 
   reg __395087_395087;
   reg _395088_395088 ; 
   reg __395088_395088;
   reg _395089_395089 ; 
   reg __395089_395089;
   reg _395090_395090 ; 
   reg __395090_395090;
   reg _395091_395091 ; 
   reg __395091_395091;
   reg _395092_395092 ; 
   reg __395092_395092;
   reg _395093_395093 ; 
   reg __395093_395093;
   reg _395094_395094 ; 
   reg __395094_395094;
   reg _395095_395095 ; 
   reg __395095_395095;
   reg _395096_395096 ; 
   reg __395096_395096;
   reg _395097_395097 ; 
   reg __395097_395097;
   reg _395098_395098 ; 
   reg __395098_395098;
   reg _395099_395099 ; 
   reg __395099_395099;
   reg _395100_395100 ; 
   reg __395100_395100;
   reg _395101_395101 ; 
   reg __395101_395101;
   reg _395102_395102 ; 
   reg __395102_395102;
   reg _395103_395103 ; 
   reg __395103_395103;
   reg _395104_395104 ; 
   reg __395104_395104;
   reg _395105_395105 ; 
   reg __395105_395105;
   reg _395106_395106 ; 
   reg __395106_395106;
   reg _395107_395107 ; 
   reg __395107_395107;
   reg _395108_395108 ; 
   reg __395108_395108;
   reg _395109_395109 ; 
   reg __395109_395109;
   reg _395110_395110 ; 
   reg __395110_395110;
   reg _395111_395111 ; 
   reg __395111_395111;
   reg _395112_395112 ; 
   reg __395112_395112;
   reg _395113_395113 ; 
   reg __395113_395113;
   reg _395114_395114 ; 
   reg __395114_395114;
   reg _395115_395115 ; 
   reg __395115_395115;
   reg _395116_395116 ; 
   reg __395116_395116;
   reg _395117_395117 ; 
   reg __395117_395117;
   reg _395118_395118 ; 
   reg __395118_395118;
   reg _395119_395119 ; 
   reg __395119_395119;
   reg _395120_395120 ; 
   reg __395120_395120;
   reg _395121_395121 ; 
   reg __395121_395121;
   reg _395122_395122 ; 
   reg __395122_395122;
   reg _395123_395123 ; 
   reg __395123_395123;
   reg _395124_395124 ; 
   reg __395124_395124;
   reg _395125_395125 ; 
   reg __395125_395125;
   reg _395126_395126 ; 
   reg __395126_395126;
   reg _395127_395127 ; 
   reg __395127_395127;
   reg _395128_395128 ; 
   reg __395128_395128;
   reg _395129_395129 ; 
   reg __395129_395129;
   reg _395130_395130 ; 
   reg __395130_395130;
   reg _395131_395131 ; 
   reg __395131_395131;
   reg _395132_395132 ; 
   reg __395132_395132;
   reg _395133_395133 ; 
   reg __395133_395133;
   reg _395134_395134 ; 
   reg __395134_395134;
   reg _395135_395135 ; 
   reg __395135_395135;
   reg _395136_395136 ; 
   reg __395136_395136;
   reg _395137_395137 ; 
   reg __395137_395137;
   reg _395138_395138 ; 
   reg __395138_395138;
   reg _395139_395139 ; 
   reg __395139_395139;
   reg _395140_395140 ; 
   reg __395140_395140;
   reg _395141_395141 ; 
   reg __395141_395141;
   reg _395142_395142 ; 
   reg __395142_395142;
   reg _395143_395143 ; 
   reg __395143_395143;
   reg _395144_395144 ; 
   reg __395144_395144;
   reg _395145_395145 ; 
   reg __395145_395145;
   reg _395146_395146 ; 
   reg __395146_395146;
   reg _395147_395147 ; 
   reg __395147_395147;
   reg _395148_395148 ; 
   reg __395148_395148;
   reg _395149_395149 ; 
   reg __395149_395149;
   reg _395150_395150 ; 
   reg __395150_395150;
   reg _395151_395151 ; 
   reg __395151_395151;
   reg _395152_395152 ; 
   reg __395152_395152;
   reg _395153_395153 ; 
   reg __395153_395153;
   reg _395154_395154 ; 
   reg __395154_395154;
   reg _395155_395155 ; 
   reg __395155_395155;
   reg _395156_395156 ; 
   reg __395156_395156;
   reg _395157_395157 ; 
   reg __395157_395157;
   reg _395158_395158 ; 
   reg __395158_395158;
   reg _395159_395159 ; 
   reg __395159_395159;
   reg _395160_395160 ; 
   reg __395160_395160;
   reg _395161_395161 ; 
   reg __395161_395161;
   reg _395162_395162 ; 
   reg __395162_395162;
   reg _395163_395163 ; 
   reg __395163_395163;
   reg _395164_395164 ; 
   reg __395164_395164;
   reg _395165_395165 ; 
   reg __395165_395165;
   reg _395166_395166 ; 
   reg __395166_395166;
   reg _395167_395167 ; 
   reg __395167_395167;
   reg _395168_395168 ; 
   reg __395168_395168;
   reg _395169_395169 ; 
   reg __395169_395169;
   reg _395170_395170 ; 
   reg __395170_395170;
   reg _395171_395171 ; 
   reg __395171_395171;
   reg _395172_395172 ; 
   reg __395172_395172;
   reg _395173_395173 ; 
   reg __395173_395173;
   reg _395174_395174 ; 
   reg __395174_395174;
   reg _395175_395175 ; 
   reg __395175_395175;
   reg _395176_395176 ; 
   reg __395176_395176;
   reg _395177_395177 ; 
   reg __395177_395177;
   reg _395178_395178 ; 
   reg __395178_395178;
   reg _395179_395179 ; 
   reg __395179_395179;
   reg _395180_395180 ; 
   reg __395180_395180;
   reg _395181_395181 ; 
   reg __395181_395181;
   reg _395182_395182 ; 
   reg __395182_395182;
   reg _395183_395183 ; 
   reg __395183_395183;
   reg _395184_395184 ; 
   reg __395184_395184;
   reg _395185_395185 ; 
   reg __395185_395185;
   reg _395186_395186 ; 
   reg __395186_395186;
   reg _395187_395187 ; 
   reg __395187_395187;
   reg _395188_395188 ; 
   reg __395188_395188;
   reg _395189_395189 ; 
   reg __395189_395189;
   reg _395190_395190 ; 
   reg __395190_395190;
   reg _395191_395191 ; 
   reg __395191_395191;
   reg _395192_395192 ; 
   reg __395192_395192;
   reg _395193_395193 ; 
   reg __395193_395193;
   reg _395194_395194 ; 
   reg __395194_395194;
   reg _395195_395195 ; 
   reg __395195_395195;
   reg _395196_395196 ; 
   reg __395196_395196;
   reg _395197_395197 ; 
   reg __395197_395197;
   reg _395198_395198 ; 
   reg __395198_395198;
   reg _395199_395199 ; 
   reg __395199_395199;
   reg _395200_395200 ; 
   reg __395200_395200;
   reg _395201_395201 ; 
   reg __395201_395201;
   reg _395202_395202 ; 
   reg __395202_395202;
   reg _395203_395203 ; 
   reg __395203_395203;
   reg _395204_395204 ; 
   reg __395204_395204;
   reg _395205_395205 ; 
   reg __395205_395205;
   reg _395206_395206 ; 
   reg __395206_395206;
   reg _395207_395207 ; 
   reg __395207_395207;
   reg _395208_395208 ; 
   reg __395208_395208;
   reg _395209_395209 ; 
   reg __395209_395209;
   reg _395210_395210 ; 
   reg __395210_395210;
   reg _395211_395211 ; 
   reg __395211_395211;
   reg _395212_395212 ; 
   reg __395212_395212;
   reg _395213_395213 ; 
   reg __395213_395213;
   reg _395214_395214 ; 
   reg __395214_395214;
   reg _395215_395215 ; 
   reg __395215_395215;
   reg _395216_395216 ; 
   reg __395216_395216;
   reg _395217_395217 ; 
   reg __395217_395217;
   reg _395218_395218 ; 
   reg __395218_395218;
   reg _395219_395219 ; 
   reg __395219_395219;
   reg _395220_395220 ; 
   reg __395220_395220;
   reg _395221_395221 ; 
   reg __395221_395221;
   reg _395222_395222 ; 
   reg __395222_395222;
   reg _395223_395223 ; 
   reg __395223_395223;
   reg _395224_395224 ; 
   reg __395224_395224;
   reg _395225_395225 ; 
   reg __395225_395225;
   reg _395226_395226 ; 
   reg __395226_395226;
   reg _395227_395227 ; 
   reg __395227_395227;
   reg _395228_395228 ; 
   reg __395228_395228;
   reg _395229_395229 ; 
   reg __395229_395229;
   reg _395230_395230 ; 
   reg __395230_395230;
   reg _395231_395231 ; 
   reg __395231_395231;
   reg _395232_395232 ; 
   reg __395232_395232;
   reg _395233_395233 ; 
   reg __395233_395233;
   reg _395234_395234 ; 
   reg __395234_395234;
   reg _395235_395235 ; 
   reg __395235_395235;
   reg _395236_395236 ; 
   reg __395236_395236;
   reg _395237_395237 ; 
   reg __395237_395237;
   reg _395238_395238 ; 
   reg __395238_395238;
   reg _395239_395239 ; 
   reg __395239_395239;
   reg _395240_395240 ; 
   reg __395240_395240;
   reg _395241_395241 ; 
   reg __395241_395241;
   reg _395242_395242 ; 
   reg __395242_395242;
   reg _395243_395243 ; 
   reg __395243_395243;
   reg _395244_395244 ; 
   reg __395244_395244;
   reg _395245_395245 ; 
   reg __395245_395245;
   reg _395246_395246 ; 
   reg __395246_395246;
   reg _395247_395247 ; 
   reg __395247_395247;
   reg _395248_395248 ; 
   reg __395248_395248;
   reg _395249_395249 ; 
   reg __395249_395249;
   reg _395250_395250 ; 
   reg __395250_395250;
   reg _395251_395251 ; 
   reg __395251_395251;
   reg _395252_395252 ; 
   reg __395252_395252;
   reg _395253_395253 ; 
   reg __395253_395253;
   reg _395254_395254 ; 
   reg __395254_395254;
   reg _395255_395255 ; 
   reg __395255_395255;
   reg _395256_395256 ; 
   reg __395256_395256;
   reg _395257_395257 ; 
   reg __395257_395257;
   reg _395258_395258 ; 
   reg __395258_395258;
   reg _395259_395259 ; 
   reg __395259_395259;
   reg _395260_395260 ; 
   reg __395260_395260;
   reg _395261_395261 ; 
   reg __395261_395261;
   reg _395262_395262 ; 
   reg __395262_395262;
   reg _395263_395263 ; 
   reg __395263_395263;
   reg _395264_395264 ; 
   reg __395264_395264;
   reg _395265_395265 ; 
   reg __395265_395265;
   reg _395266_395266 ; 
   reg __395266_395266;
   reg _395267_395267 ; 
   reg __395267_395267;
   reg _395268_395268 ; 
   reg __395268_395268;
   reg _395269_395269 ; 
   reg __395269_395269;
   reg _395270_395270 ; 
   reg __395270_395270;
   reg _395271_395271 ; 
   reg __395271_395271;
   reg _395272_395272 ; 
   reg __395272_395272;
   reg _395273_395273 ; 
   reg __395273_395273;
   reg _395274_395274 ; 
   reg __395274_395274;
   reg _395275_395275 ; 
   reg __395275_395275;
   reg _395276_395276 ; 
   reg __395276_395276;
   reg _395277_395277 ; 
   reg __395277_395277;
   reg _395278_395278 ; 
   reg __395278_395278;
   reg _395279_395279 ; 
   reg __395279_395279;
   reg _395280_395280 ; 
   reg __395280_395280;
   reg _395281_395281 ; 
   reg __395281_395281;
   reg _395282_395282 ; 
   reg __395282_395282;
   reg _395283_395283 ; 
   reg __395283_395283;
   reg _395284_395284 ; 
   reg __395284_395284;
   reg _395285_395285 ; 
   reg __395285_395285;
   reg _395286_395286 ; 
   reg __395286_395286;
   reg _395287_395287 ; 
   reg __395287_395287;
   reg _395288_395288 ; 
   reg __395288_395288;
   reg _395289_395289 ; 
   reg __395289_395289;
   reg _395290_395290 ; 
   reg __395290_395290;
   reg _395291_395291 ; 
   reg __395291_395291;
   reg _395292_395292 ; 
   reg __395292_395292;
   reg _395293_395293 ; 
   reg __395293_395293;
   reg _395294_395294 ; 
   reg __395294_395294;
   reg _395295_395295 ; 
   reg __395295_395295;
   reg _395296_395296 ; 
   reg __395296_395296;
   reg _395297_395297 ; 
   reg __395297_395297;
   reg _395298_395298 ; 
   reg __395298_395298;
   reg _395299_395299 ; 
   reg __395299_395299;
   reg _395300_395300 ; 
   reg __395300_395300;
   reg _395301_395301 ; 
   reg __395301_395301;
   reg _395302_395302 ; 
   reg __395302_395302;
   reg _395303_395303 ; 
   reg __395303_395303;
   reg _395304_395304 ; 
   reg __395304_395304;
   reg _395305_395305 ; 
   reg __395305_395305;
   reg _395306_395306 ; 
   reg __395306_395306;
   reg _395307_395307 ; 
   reg __395307_395307;
   reg _395308_395308 ; 
   reg __395308_395308;
   reg _395309_395309 ; 
   reg __395309_395309;
   reg _395310_395310 ; 
   reg __395310_395310;
   reg _395311_395311 ; 
   reg __395311_395311;
   reg _395312_395312 ; 
   reg __395312_395312;
   reg _395313_395313 ; 
   reg __395313_395313;
   reg _395314_395314 ; 
   reg __395314_395314;
   reg _395315_395315 ; 
   reg __395315_395315;
   reg _395316_395316 ; 
   reg __395316_395316;
   reg _395317_395317 ; 
   reg __395317_395317;
   reg _395318_395318 ; 
   reg __395318_395318;
   reg _395319_395319 ; 
   reg __395319_395319;
   reg _395320_395320 ; 
   reg __395320_395320;
   reg _395321_395321 ; 
   reg __395321_395321;
   reg _395322_395322 ; 
   reg __395322_395322;
   reg _395323_395323 ; 
   reg __395323_395323;
   reg _395324_395324 ; 
   reg __395324_395324;
   reg _395325_395325 ; 
   reg __395325_395325;
   reg _395326_395326 ; 
   reg __395326_395326;
   reg _395327_395327 ; 
   reg __395327_395327;
   reg _395328_395328 ; 
   reg __395328_395328;
   reg _395329_395329 ; 
   reg __395329_395329;
   reg _395330_395330 ; 
   reg __395330_395330;
   reg _395331_395331 ; 
   reg __395331_395331;
   reg _395332_395332 ; 
   reg __395332_395332;
   reg _395333_395333 ; 
   reg __395333_395333;
   reg _395334_395334 ; 
   reg __395334_395334;
   reg _395335_395335 ; 
   reg __395335_395335;
   reg _395336_395336 ; 
   reg __395336_395336;
   reg _395337_395337 ; 
   reg __395337_395337;
   reg _395338_395338 ; 
   reg __395338_395338;
   reg _395339_395339 ; 
   reg __395339_395339;
   reg _395340_395340 ; 
   reg __395340_395340;
   reg _395341_395341 ; 
   reg __395341_395341;
   reg _395342_395342 ; 
   reg __395342_395342;
   reg _395343_395343 ; 
   reg __395343_395343;
   reg _395344_395344 ; 
   reg __395344_395344;
   reg _395345_395345 ; 
   reg __395345_395345;
   reg _395346_395346 ; 
   reg __395346_395346;
   reg _395347_395347 ; 
   reg __395347_395347;
   reg _395348_395348 ; 
   reg __395348_395348;
   reg _395349_395349 ; 
   reg __395349_395349;
   reg _395350_395350 ; 
   reg __395350_395350;
   reg _395351_395351 ; 
   reg __395351_395351;
   reg _395352_395352 ; 
   reg __395352_395352;
   reg _395353_395353 ; 
   reg __395353_395353;
   reg _395354_395354 ; 
   reg __395354_395354;
   reg _395355_395355 ; 
   reg __395355_395355;
   reg _395356_395356 ; 
   reg __395356_395356;
   reg _395357_395357 ; 
   reg __395357_395357;
   reg _395358_395358 ; 
   reg __395358_395358;
   reg _395359_395359 ; 
   reg __395359_395359;
   reg _395360_395360 ; 
   reg __395360_395360;
   reg _395361_395361 ; 
   reg __395361_395361;
   reg _395362_395362 ; 
   reg __395362_395362;
   reg _395363_395363 ; 
   reg __395363_395363;
   reg _395364_395364 ; 
   reg __395364_395364;
   reg _395365_395365 ; 
   reg __395365_395365;
   reg _395366_395366 ; 
   reg __395366_395366;
   reg _395367_395367 ; 
   reg __395367_395367;
   reg _395368_395368 ; 
   reg __395368_395368;
   reg _395369_395369 ; 
   reg __395369_395369;
   reg _395370_395370 ; 
   reg __395370_395370;
   reg _395371_395371 ; 
   reg __395371_395371;
   reg _395372_395372 ; 
   reg __395372_395372;
   reg _395373_395373 ; 
   reg __395373_395373;
   reg _395374_395374 ; 
   reg __395374_395374;
   reg _395375_395375 ; 
   reg __395375_395375;
   reg _395376_395376 ; 
   reg __395376_395376;
   reg _395377_395377 ; 
   reg __395377_395377;
   reg _395378_395378 ; 
   reg __395378_395378;
   reg _395379_395379 ; 
   reg __395379_395379;
   reg _395380_395380 ; 
   reg __395380_395380;
   reg _395381_395381 ; 
   reg __395381_395381;
   reg _395382_395382 ; 
   reg __395382_395382;
   reg _395383_395383 ; 
   reg __395383_395383;
   reg _395384_395384 ; 
   reg __395384_395384;
   reg _395385_395385 ; 
   reg __395385_395385;
   reg _395386_395386 ; 
   reg __395386_395386;
   reg _395387_395387 ; 
   reg __395387_395387;
   reg _395388_395388 ; 
   reg __395388_395388;
   reg _395389_395389 ; 
   reg __395389_395389;
   reg _395390_395390 ; 
   reg __395390_395390;
   reg _395391_395391 ; 
   reg __395391_395391;
   reg _395392_395392 ; 
   reg __395392_395392;
   reg _395393_395393 ; 
   reg __395393_395393;
   reg _395394_395394 ; 
   reg __395394_395394;
   reg _395395_395395 ; 
   reg __395395_395395;
   reg _395396_395396 ; 
   reg __395396_395396;
   reg _395397_395397 ; 
   reg __395397_395397;
   reg _395398_395398 ; 
   reg __395398_395398;
   reg _395399_395399 ; 
   reg __395399_395399;
   reg _395400_395400 ; 
   reg __395400_395400;
   reg _395401_395401 ; 
   reg __395401_395401;
   reg _395402_395402 ; 
   reg __395402_395402;
   reg _395403_395403 ; 
   reg __395403_395403;
   reg _395404_395404 ; 
   reg __395404_395404;
   reg _395405_395405 ; 
   reg __395405_395405;
   reg _395406_395406 ; 
   reg __395406_395406;
   reg _395407_395407 ; 
   reg __395407_395407;
   reg _395408_395408 ; 
   reg __395408_395408;
   reg _395409_395409 ; 
   reg __395409_395409;
   reg _395410_395410 ; 
   reg __395410_395410;
   reg _395411_395411 ; 
   reg __395411_395411;
   reg _395412_395412 ; 
   reg __395412_395412;
   reg _395413_395413 ; 
   reg __395413_395413;
   reg _395414_395414 ; 
   reg __395414_395414;
   reg _395415_395415 ; 
   reg __395415_395415;
   reg _395416_395416 ; 
   reg __395416_395416;
   reg _395417_395417 ; 
   reg __395417_395417;
   reg _395418_395418 ; 
   reg __395418_395418;
   reg _395419_395419 ; 
   reg __395419_395419;
   reg _395420_395420 ; 
   reg __395420_395420;
   reg _395421_395421 ; 
   reg __395421_395421;
   reg _395422_395422 ; 
   reg __395422_395422;
   reg _395423_395423 ; 
   reg __395423_395423;
   reg _395424_395424 ; 
   reg __395424_395424;
   reg _395425_395425 ; 
   reg __395425_395425;
   reg _395426_395426 ; 
   reg __395426_395426;
   reg _395427_395427 ; 
   reg __395427_395427;
   reg _395428_395428 ; 
   reg __395428_395428;
   reg _395429_395429 ; 
   reg __395429_395429;
   reg _395430_395430 ; 
   reg __395430_395430;
   reg _395431_395431 ; 
   reg __395431_395431;
   reg _395432_395432 ; 
   reg __395432_395432;
   reg _395433_395433 ; 
   reg __395433_395433;
   reg _395434_395434 ; 
   reg __395434_395434;
   reg _395435_395435 ; 
   reg __395435_395435;
   reg _395436_395436 ; 
   reg __395436_395436;
   reg _395437_395437 ; 
   reg __395437_395437;
   reg _395438_395438 ; 
   reg __395438_395438;
   reg _395439_395439 ; 
   reg __395439_395439;
   reg _395440_395440 ; 
   reg __395440_395440;
   reg _395441_395441 ; 
   reg __395441_395441;
   reg _395442_395442 ; 
   reg __395442_395442;
   reg _395443_395443 ; 
   reg __395443_395443;
   reg _395444_395444 ; 
   reg __395444_395444;
   reg _395445_395445 ; 
   reg __395445_395445;
   reg _395446_395446 ; 
   reg __395446_395446;
   reg _395447_395447 ; 
   reg __395447_395447;
   reg _395448_395448 ; 
   reg __395448_395448;
   reg _395449_395449 ; 
   reg __395449_395449;
   reg _395450_395450 ; 
   reg __395450_395450;
   reg _395451_395451 ; 
   reg __395451_395451;
   reg _395452_395452 ; 
   reg __395452_395452;
   reg _395453_395453 ; 
   reg __395453_395453;
   reg _395454_395454 ; 
   reg __395454_395454;
   reg _395455_395455 ; 
   reg __395455_395455;
   reg _395456_395456 ; 
   reg __395456_395456;
   reg _395457_395457 ; 
   reg __395457_395457;
   reg _395458_395458 ; 
   reg __395458_395458;
   reg _395459_395459 ; 
   reg __395459_395459;
   reg _395460_395460 ; 
   reg __395460_395460;
   reg _395461_395461 ; 
   reg __395461_395461;
   reg _395462_395462 ; 
   reg __395462_395462;
   reg _395463_395463 ; 
   reg __395463_395463;
   reg _395464_395464 ; 
   reg __395464_395464;
   reg _395465_395465 ; 
   reg __395465_395465;
   reg _395466_395466 ; 
   reg __395466_395466;
   reg _395467_395467 ; 
   reg __395467_395467;
   reg _395468_395468 ; 
   reg __395468_395468;
   reg _395469_395469 ; 
   reg __395469_395469;
   reg _395470_395470 ; 
   reg __395470_395470;
   reg _395471_395471 ; 
   reg __395471_395471;
   reg _395472_395472 ; 
   reg __395472_395472;
   reg _395473_395473 ; 
   reg __395473_395473;
   reg _395474_395474 ; 
   reg __395474_395474;
   reg _395475_395475 ; 
   reg __395475_395475;
   reg _395476_395476 ; 
   reg __395476_395476;
   reg _395477_395477 ; 
   reg __395477_395477;
   reg _395478_395478 ; 
   reg __395478_395478;
   reg _395479_395479 ; 
   reg __395479_395479;
   reg _395480_395480 ; 
   reg __395480_395480;
   reg _395481_395481 ; 
   reg __395481_395481;
   reg _395482_395482 ; 
   reg __395482_395482;
   reg _395483_395483 ; 
   reg __395483_395483;
   reg _395484_395484 ; 
   reg __395484_395484;
   reg _395485_395485 ; 
   reg __395485_395485;
   reg _395486_395486 ; 
   reg __395486_395486;
   reg _395487_395487 ; 
   reg __395487_395487;
   reg _395488_395488 ; 
   reg __395488_395488;
   reg _395489_395489 ; 
   reg __395489_395489;
   reg _395490_395490 ; 
   reg __395490_395490;
   reg _395491_395491 ; 
   reg __395491_395491;
   reg _395492_395492 ; 
   reg __395492_395492;
   reg _395493_395493 ; 
   reg __395493_395493;
   reg _395494_395494 ; 
   reg __395494_395494;
   reg _395495_395495 ; 
   reg __395495_395495;
   reg _395496_395496 ; 
   reg __395496_395496;
   reg _395497_395497 ; 
   reg __395497_395497;
   reg _395498_395498 ; 
   reg __395498_395498;
   reg _395499_395499 ; 
   reg __395499_395499;
   reg _395500_395500 ; 
   reg __395500_395500;
   reg _395501_395501 ; 
   reg __395501_395501;
   reg _395502_395502 ; 
   reg __395502_395502;
   reg _395503_395503 ; 
   reg __395503_395503;
   reg _395504_395504 ; 
   reg __395504_395504;
   reg _395505_395505 ; 
   reg __395505_395505;
   reg _395506_395506 ; 
   reg __395506_395506;
   reg _395507_395507 ; 
   reg __395507_395507;
   reg _395508_395508 ; 
   reg __395508_395508;
   reg _395509_395509 ; 
   reg __395509_395509;
   reg _395510_395510 ; 
   reg __395510_395510;
   reg _395511_395511 ; 
   reg __395511_395511;
   reg _395512_395512 ; 
   reg __395512_395512;
   reg _395513_395513 ; 
   reg __395513_395513;
   reg _395514_395514 ; 
   reg __395514_395514;
   reg _395515_395515 ; 
   reg __395515_395515;
   reg _395516_395516 ; 
   reg __395516_395516;
   reg _395517_395517 ; 
   reg __395517_395517;
   reg _395518_395518 ; 
   reg __395518_395518;
   reg _395519_395519 ; 
   reg __395519_395519;
   reg _395520_395520 ; 
   reg __395520_395520;
   reg _395521_395521 ; 
   reg __395521_395521;
   reg _395522_395522 ; 
   reg __395522_395522;
   reg _395523_395523 ; 
   reg __395523_395523;
   reg _395524_395524 ; 
   reg __395524_395524;
   reg _395525_395525 ; 
   reg __395525_395525;
   reg _395526_395526 ; 
   reg __395526_395526;
   reg _395527_395527 ; 
   reg __395527_395527;
   reg _395528_395528 ; 
   reg __395528_395528;
   reg _395529_395529 ; 
   reg __395529_395529;
   reg _395530_395530 ; 
   reg __395530_395530;
   reg _395531_395531 ; 
   reg __395531_395531;
   reg _395532_395532 ; 
   reg __395532_395532;
   reg _395533_395533 ; 
   reg __395533_395533;
   reg _395534_395534 ; 
   reg __395534_395534;
   reg _395535_395535 ; 
   reg __395535_395535;
   reg _395536_395536 ; 
   reg __395536_395536;
   reg _395537_395537 ; 
   reg __395537_395537;
   reg _395538_395538 ; 
   reg __395538_395538;
   reg _395539_395539 ; 
   reg __395539_395539;
   reg _395540_395540 ; 
   reg __395540_395540;
   reg _395541_395541 ; 
   reg __395541_395541;
   reg _395542_395542 ; 
   reg __395542_395542;
   reg _395543_395543 ; 
   reg __395543_395543;
   reg _395544_395544 ; 
   reg __395544_395544;
   reg _395545_395545 ; 
   reg __395545_395545;
   reg _395546_395546 ; 
   reg __395546_395546;
   reg _395547_395547 ; 
   reg __395547_395547;
   reg _395548_395548 ; 
   reg __395548_395548;
   reg _395549_395549 ; 
   reg __395549_395549;
   reg _395550_395550 ; 
   reg __395550_395550;
   reg _395551_395551 ; 
   reg __395551_395551;
   reg _395552_395552 ; 
   reg __395552_395552;
   reg _395553_395553 ; 
   reg __395553_395553;
   reg _395554_395554 ; 
   reg __395554_395554;
   reg _395555_395555 ; 
   reg __395555_395555;
   reg _395556_395556 ; 
   reg __395556_395556;
   reg _395557_395557 ; 
   reg __395557_395557;
   reg _395558_395558 ; 
   reg __395558_395558;
   reg _395559_395559 ; 
   reg __395559_395559;
   reg _395560_395560 ; 
   reg __395560_395560;
   reg _395561_395561 ; 
   reg __395561_395561;
   reg _395562_395562 ; 
   reg __395562_395562;
   reg _395563_395563 ; 
   reg __395563_395563;
   reg _395564_395564 ; 
   reg __395564_395564;
   reg _395565_395565 ; 
   reg __395565_395565;
   reg _395566_395566 ; 
   reg __395566_395566;
   reg _395567_395567 ; 
   reg __395567_395567;
   reg _395568_395568 ; 
   reg __395568_395568;
   reg _395569_395569 ; 
   reg __395569_395569;
   reg _395570_395570 ; 
   reg __395570_395570;
   reg _395571_395571 ; 
   reg __395571_395571;
   reg _395572_395572 ; 
   reg __395572_395572;
   reg _395573_395573 ; 
   reg __395573_395573;
   reg _395574_395574 ; 
   reg __395574_395574;
   reg _395575_395575 ; 
   reg __395575_395575;
   reg _395576_395576 ; 
   reg __395576_395576;
   reg _395577_395577 ; 
   reg __395577_395577;
   reg _395578_395578 ; 
   reg __395578_395578;
   reg _395579_395579 ; 
   reg __395579_395579;
   reg _395580_395580 ; 
   reg __395580_395580;
   reg _395581_395581 ; 
   reg __395581_395581;
   reg _395582_395582 ; 
   reg __395582_395582;
   reg _395583_395583 ; 
   reg __395583_395583;
   reg _395584_395584 ; 
   reg __395584_395584;
   reg _395585_395585 ; 
   reg __395585_395585;
   reg _395586_395586 ; 
   reg __395586_395586;
   reg _395587_395587 ; 
   reg __395587_395587;
   reg _395588_395588 ; 
   reg __395588_395588;
   reg _395589_395589 ; 
   reg __395589_395589;
   reg _395590_395590 ; 
   reg __395590_395590;
   reg _395591_395591 ; 
   reg __395591_395591;
   reg _395592_395592 ; 
   reg __395592_395592;
   reg _395593_395593 ; 
   reg __395593_395593;
   reg _395594_395594 ; 
   reg __395594_395594;
   reg _395595_395595 ; 
   reg __395595_395595;
   reg _395596_395596 ; 
   reg __395596_395596;
   reg _395597_395597 ; 
   reg __395597_395597;
   reg _395598_395598 ; 
   reg __395598_395598;
   reg _395599_395599 ; 
   reg __395599_395599;
   reg _395600_395600 ; 
   reg __395600_395600;
   reg _395601_395601 ; 
   reg __395601_395601;
   reg _395602_395602 ; 
   reg __395602_395602;
   reg _395603_395603 ; 
   reg __395603_395603;
   reg _395604_395604 ; 
   reg __395604_395604;
   reg _395605_395605 ; 
   reg __395605_395605;
   reg _395606_395606 ; 
   reg __395606_395606;
   reg _395607_395607 ; 
   reg __395607_395607;
   reg _395608_395608 ; 
   reg __395608_395608;
   reg _395609_395609 ; 
   reg __395609_395609;
   reg _395610_395610 ; 
   reg __395610_395610;
   reg _395611_395611 ; 
   reg __395611_395611;
   reg _395612_395612 ; 
   reg __395612_395612;
   reg _395613_395613 ; 
   reg __395613_395613;
   reg _395614_395614 ; 
   reg __395614_395614;
   reg _395615_395615 ; 
   reg __395615_395615;
   reg _395616_395616 ; 
   reg __395616_395616;
   reg _395617_395617 ; 
   reg __395617_395617;
   reg _395618_395618 ; 
   reg __395618_395618;
   reg _395619_395619 ; 
   reg __395619_395619;
   reg _395620_395620 ; 
   reg __395620_395620;
   reg _395621_395621 ; 
   reg __395621_395621;
   reg _395622_395622 ; 
   reg __395622_395622;
   reg _395623_395623 ; 
   reg __395623_395623;
   reg _395624_395624 ; 
   reg __395624_395624;
   reg _395625_395625 ; 
   reg __395625_395625;
   reg _395626_395626 ; 
   reg __395626_395626;
   reg _395627_395627 ; 
   reg __395627_395627;
   reg _395628_395628 ; 
   reg __395628_395628;
   reg _395629_395629 ; 
   reg __395629_395629;
   reg _395630_395630 ; 
   reg __395630_395630;
   reg _395631_395631 ; 
   reg __395631_395631;
   reg _395632_395632 ; 
   reg __395632_395632;
   reg _395633_395633 ; 
   reg __395633_395633;
   reg _395634_395634 ; 
   reg __395634_395634;
   reg _395635_395635 ; 
   reg __395635_395635;
   reg _395636_395636 ; 
   reg __395636_395636;
   reg _395637_395637 ; 
   reg __395637_395637;
   reg _395638_395638 ; 
   reg __395638_395638;
   reg _395639_395639 ; 
   reg __395639_395639;
   reg _395640_395640 ; 
   reg __395640_395640;
   reg _395641_395641 ; 
   reg __395641_395641;
   reg _395642_395642 ; 
   reg __395642_395642;
   reg _395643_395643 ; 
   reg __395643_395643;
   reg _395644_395644 ; 
   reg __395644_395644;
   reg _395645_395645 ; 
   reg __395645_395645;
   reg _395646_395646 ; 
   reg __395646_395646;
   reg _395647_395647 ; 
   reg __395647_395647;
   reg _395648_395648 ; 
   reg __395648_395648;
   reg _395649_395649 ; 
   reg __395649_395649;
   reg _395650_395650 ; 
   reg __395650_395650;
   reg _395651_395651 ; 
   reg __395651_395651;
   reg _395652_395652 ; 
   reg __395652_395652;
   reg _395653_395653 ; 
   reg __395653_395653;
   reg _395654_395654 ; 
   reg __395654_395654;
   reg _395655_395655 ; 
   reg __395655_395655;
   reg _395656_395656 ; 
   reg __395656_395656;
   reg _395657_395657 ; 
   reg __395657_395657;
   reg _395658_395658 ; 
   reg __395658_395658;
   reg _395659_395659 ; 
   reg __395659_395659;
   reg _395660_395660 ; 
   reg __395660_395660;
   reg _395661_395661 ; 
   reg __395661_395661;
   reg _395662_395662 ; 
   reg __395662_395662;
   reg _395663_395663 ; 
   reg __395663_395663;
   reg _395664_395664 ; 
   reg __395664_395664;
   reg _395665_395665 ; 
   reg __395665_395665;
   reg _395666_395666 ; 
   reg __395666_395666;
   reg _395667_395667 ; 
   reg __395667_395667;
   reg _395668_395668 ; 
   reg __395668_395668;
   reg _395669_395669 ; 
   reg __395669_395669;
   reg _395670_395670 ; 
   reg __395670_395670;
   reg _395671_395671 ; 
   reg __395671_395671;
   reg _395672_395672 ; 
   reg __395672_395672;
   reg _395673_395673 ; 
   reg __395673_395673;
   reg _395674_395674 ; 
   reg __395674_395674;
   reg _395675_395675 ; 
   reg __395675_395675;
   reg _395676_395676 ; 
   reg __395676_395676;
   reg _395677_395677 ; 
   reg __395677_395677;
   reg _395678_395678 ; 
   reg __395678_395678;
   reg _395679_395679 ; 
   reg __395679_395679;
   reg _395680_395680 ; 
   reg __395680_395680;
   reg _395681_395681 ; 
   reg __395681_395681;
   reg _395682_395682 ; 
   reg __395682_395682;
   reg _395683_395683 ; 
   reg __395683_395683;
   reg _395684_395684 ; 
   reg __395684_395684;
   reg _395685_395685 ; 
   reg __395685_395685;
   reg _395686_395686 ; 
   reg __395686_395686;
   reg _395687_395687 ; 
   reg __395687_395687;
   reg _395688_395688 ; 
   reg __395688_395688;
   reg _395689_395689 ; 
   reg __395689_395689;
   reg _395690_395690 ; 
   reg __395690_395690;
   reg _395691_395691 ; 
   reg __395691_395691;
   reg _395692_395692 ; 
   reg __395692_395692;
   reg _395693_395693 ; 
   reg __395693_395693;
   reg _395694_395694 ; 
   reg __395694_395694;
   reg _395695_395695 ; 
   reg __395695_395695;
   reg _395696_395696 ; 
   reg __395696_395696;
   reg _395697_395697 ; 
   reg __395697_395697;
   reg _395698_395698 ; 
   reg __395698_395698;
   reg _395699_395699 ; 
   reg __395699_395699;
   reg _395700_395700 ; 
   reg __395700_395700;
   reg _395701_395701 ; 
   reg __395701_395701;
   reg _395702_395702 ; 
   reg __395702_395702;
   reg _395703_395703 ; 
   reg __395703_395703;
   reg _395704_395704 ; 
   reg __395704_395704;
   reg _395705_395705 ; 
   reg __395705_395705;
   reg _395706_395706 ; 
   reg __395706_395706;
   reg _395707_395707 ; 
   reg __395707_395707;
   reg _395708_395708 ; 
   reg __395708_395708;
   reg _395709_395709 ; 
   reg __395709_395709;
   reg _395710_395710 ; 
   reg __395710_395710;
   reg _395711_395711 ; 
   reg __395711_395711;
   reg _395712_395712 ; 
   reg __395712_395712;
   reg _395713_395713 ; 
   reg __395713_395713;
   reg _395714_395714 ; 
   reg __395714_395714;
   reg _395715_395715 ; 
   reg __395715_395715;
   reg _395716_395716 ; 
   reg __395716_395716;
   reg _395717_395717 ; 
   reg __395717_395717;
   reg _395718_395718 ; 
   reg __395718_395718;
   reg _395719_395719 ; 
   reg __395719_395719;
   reg _395720_395720 ; 
   reg __395720_395720;
   reg _395721_395721 ; 
   reg __395721_395721;
   reg _395722_395722 ; 
   reg __395722_395722;
   reg _395723_395723 ; 
   reg __395723_395723;
   reg _395724_395724 ; 
   reg __395724_395724;
   reg _395725_395725 ; 
   reg __395725_395725;
   reg _395726_395726 ; 
   reg __395726_395726;
   reg _395727_395727 ; 
   reg __395727_395727;
   reg _395728_395728 ; 
   reg __395728_395728;
   reg _395729_395729 ; 
   reg __395729_395729;
   reg _395730_395730 ; 
   reg __395730_395730;
   reg _395731_395731 ; 
   reg __395731_395731;
   reg _395732_395732 ; 
   reg __395732_395732;
   reg _395733_395733 ; 
   reg __395733_395733;
   reg _395734_395734 ; 
   reg __395734_395734;
   reg _395735_395735 ; 
   reg __395735_395735;
   reg _395736_395736 ; 
   reg __395736_395736;
   reg _395737_395737 ; 
   reg __395737_395737;
   reg _395738_395738 ; 
   reg __395738_395738;
   reg _395739_395739 ; 
   reg __395739_395739;
   reg _395740_395740 ; 
   reg __395740_395740;
   reg _395741_395741 ; 
   reg __395741_395741;
   reg _395742_395742 ; 
   reg __395742_395742;
   reg _395743_395743 ; 
   reg __395743_395743;
   reg _395744_395744 ; 
   reg __395744_395744;
   reg _395745_395745 ; 
   reg __395745_395745;
   reg _395746_395746 ; 
   reg __395746_395746;
   reg _395747_395747 ; 
   reg __395747_395747;
   reg _395748_395748 ; 
   reg __395748_395748;
   reg _395749_395749 ; 
   reg __395749_395749;
   reg _395750_395750 ; 
   reg __395750_395750;
   reg _395751_395751 ; 
   reg __395751_395751;
   reg _395752_395752 ; 
   reg __395752_395752;
   reg _395753_395753 ; 
   reg __395753_395753;
   reg _395754_395754 ; 
   reg __395754_395754;
   reg _395755_395755 ; 
   reg __395755_395755;
   reg _395756_395756 ; 
   reg __395756_395756;
   reg _395757_395757 ; 
   reg __395757_395757;
   reg _395758_395758 ; 
   reg __395758_395758;
   reg _395759_395759 ; 
   reg __395759_395759;
   reg _395760_395760 ; 
   reg __395760_395760;
   reg _395761_395761 ; 
   reg __395761_395761;
   reg _395762_395762 ; 
   reg __395762_395762;
   reg _395763_395763 ; 
   reg __395763_395763;
   reg _395764_395764 ; 
   reg __395764_395764;
   reg _395765_395765 ; 
   reg __395765_395765;
   reg _395766_395766 ; 
   reg __395766_395766;
   reg _395767_395767 ; 
   reg __395767_395767;
   reg _395768_395768 ; 
   reg __395768_395768;
   reg _395769_395769 ; 
   reg __395769_395769;
   reg _395770_395770 ; 
   reg __395770_395770;
   reg _395771_395771 ; 
   reg __395771_395771;
   reg _395772_395772 ; 
   reg __395772_395772;
   reg _395773_395773 ; 
   reg __395773_395773;
   reg _395774_395774 ; 
   reg __395774_395774;
   reg _395775_395775 ; 
   reg __395775_395775;
   reg _395776_395776 ; 
   reg __395776_395776;
   reg _395777_395777 ; 
   reg __395777_395777;
   reg _395778_395778 ; 
   reg __395778_395778;
   reg _395779_395779 ; 
   reg __395779_395779;
   reg _395780_395780 ; 
   reg __395780_395780;
   reg _395781_395781 ; 
   reg __395781_395781;
   reg _395782_395782 ; 
   reg __395782_395782;
   reg _395783_395783 ; 
   reg __395783_395783;
   reg _395784_395784 ; 
   reg __395784_395784;
   reg _395785_395785 ; 
   reg __395785_395785;
   reg _395786_395786 ; 
   reg __395786_395786;
   reg _395787_395787 ; 
   reg __395787_395787;
   reg _395788_395788 ; 
   reg __395788_395788;
   reg _395789_395789 ; 
   reg __395789_395789;
   reg _395790_395790 ; 
   reg __395790_395790;
   reg _395791_395791 ; 
   reg __395791_395791;
   reg _395792_395792 ; 
   reg __395792_395792;
   reg _395793_395793 ; 
   reg __395793_395793;
   reg _395794_395794 ; 
   reg __395794_395794;
   reg _395795_395795 ; 
   reg __395795_395795;
   reg _395796_395796 ; 
   reg __395796_395796;
   reg _395797_395797 ; 
   reg __395797_395797;
   reg _395798_395798 ; 
   reg __395798_395798;
   reg _395799_395799 ; 
   reg __395799_395799;
   reg _395800_395800 ; 
   reg __395800_395800;
   reg _395801_395801 ; 
   reg __395801_395801;
   reg _395802_395802 ; 
   reg __395802_395802;
   reg _395803_395803 ; 
   reg __395803_395803;
   reg _395804_395804 ; 
   reg __395804_395804;
   reg _395805_395805 ; 
   reg __395805_395805;
   reg _395806_395806 ; 
   reg __395806_395806;
   reg _395807_395807 ; 
   reg __395807_395807;
   reg _395808_395808 ; 
   reg __395808_395808;
   reg _395809_395809 ; 
   reg __395809_395809;
   reg _395810_395810 ; 
   reg __395810_395810;
   reg _395811_395811 ; 
   reg __395811_395811;
   reg _395812_395812 ; 
   reg __395812_395812;
   reg _395813_395813 ; 
   reg __395813_395813;
   reg _395814_395814 ; 
   reg __395814_395814;
   reg _395815_395815 ; 
   reg __395815_395815;
   reg _395816_395816 ; 
   reg __395816_395816;
   reg _395817_395817 ; 
   reg __395817_395817;
   reg _395818_395818 ; 
   reg __395818_395818;
   reg _395819_395819 ; 
   reg __395819_395819;
   reg _395820_395820 ; 
   reg __395820_395820;
   reg _395821_395821 ; 
   reg __395821_395821;
   reg _395822_395822 ; 
   reg __395822_395822;
   reg _395823_395823 ; 
   reg __395823_395823;
   reg _395824_395824 ; 
   reg __395824_395824;
   reg _395825_395825 ; 
   reg __395825_395825;
   reg _395826_395826 ; 
   reg __395826_395826;
   reg _395827_395827 ; 
   reg __395827_395827;
   reg _395828_395828 ; 
   reg __395828_395828;
   reg _395829_395829 ; 
   reg __395829_395829;
   reg _395830_395830 ; 
   reg __395830_395830;
   reg _395831_395831 ; 
   reg __395831_395831;
   reg _395832_395832 ; 
   reg __395832_395832;
   reg _395833_395833 ; 
   reg __395833_395833;
   reg _395834_395834 ; 
   reg __395834_395834;
   reg _395835_395835 ; 
   reg __395835_395835;
   reg _395836_395836 ; 
   reg __395836_395836;
   reg _395837_395837 ; 
   reg __395837_395837;
   reg _395838_395838 ; 
   reg __395838_395838;
   reg _395839_395839 ; 
   reg __395839_395839;
   reg _395840_395840 ; 
   reg __395840_395840;
   reg _395841_395841 ; 
   reg __395841_395841;
   reg _395842_395842 ; 
   reg __395842_395842;
   reg _395843_395843 ; 
   reg __395843_395843;
   reg _395844_395844 ; 
   reg __395844_395844;
   reg _395845_395845 ; 
   reg __395845_395845;
   reg _395846_395846 ; 
   reg __395846_395846;
   reg _395847_395847 ; 
   reg __395847_395847;
   reg _395848_395848 ; 
   reg __395848_395848;
   reg _395849_395849 ; 
   reg __395849_395849;
   reg _395850_395850 ; 
   reg __395850_395850;
   reg _395851_395851 ; 
   reg __395851_395851;
   reg _395852_395852 ; 
   reg __395852_395852;
   reg _395853_395853 ; 
   reg __395853_395853;
   reg _395854_395854 ; 
   reg __395854_395854;
   reg _395855_395855 ; 
   reg __395855_395855;
   reg _395856_395856 ; 
   reg __395856_395856;
   reg _395857_395857 ; 
   reg __395857_395857;
   reg _395858_395858 ; 
   reg __395858_395858;
   reg _395859_395859 ; 
   reg __395859_395859;
   reg _395860_395860 ; 
   reg __395860_395860;
   reg _395861_395861 ; 
   reg __395861_395861;
   reg _395862_395862 ; 
   reg __395862_395862;
   reg _395863_395863 ; 
   reg __395863_395863;
   reg _395864_395864 ; 
   reg __395864_395864;
   reg _395865_395865 ; 
   reg __395865_395865;
   reg _395866_395866 ; 
   reg __395866_395866;
   reg _395867_395867 ; 
   reg __395867_395867;
   reg _395868_395868 ; 
   reg __395868_395868;
   reg _395869_395869 ; 
   reg __395869_395869;
   reg _395870_395870 ; 
   reg __395870_395870;
   reg _395871_395871 ; 
   reg __395871_395871;
   reg _395872_395872 ; 
   reg __395872_395872;
   reg _395873_395873 ; 
   reg __395873_395873;
   reg _395874_395874 ; 
   reg __395874_395874;
   reg _395875_395875 ; 
   reg __395875_395875;
   reg _395876_395876 ; 
   reg __395876_395876;
   reg _395877_395877 ; 
   reg __395877_395877;
   reg _395878_395878 ; 
   reg __395878_395878;
   reg _395879_395879 ; 
   reg __395879_395879;
   reg _395880_395880 ; 
   reg __395880_395880;
   reg _395881_395881 ; 
   reg __395881_395881;
   reg _395882_395882 ; 
   reg __395882_395882;
   reg _395883_395883 ; 
   reg __395883_395883;
   reg _395884_395884 ; 
   reg __395884_395884;
   reg _395885_395885 ; 
   reg __395885_395885;
   reg _395886_395886 ; 
   reg __395886_395886;
   reg _395887_395887 ; 
   reg __395887_395887;
   reg _395888_395888 ; 
   reg __395888_395888;
   reg _395889_395889 ; 
   reg __395889_395889;
   reg _395890_395890 ; 
   reg __395890_395890;
   reg _395891_395891 ; 
   reg __395891_395891;
   reg _395892_395892 ; 
   reg __395892_395892;
   reg _395893_395893 ; 
   reg __395893_395893;
   reg _395894_395894 ; 
   reg __395894_395894;
   reg _395895_395895 ; 
   reg __395895_395895;
   reg _395896_395896 ; 
   reg __395896_395896;
   reg _395897_395897 ; 
   reg __395897_395897;
   reg _395898_395898 ; 
   reg __395898_395898;
   reg _395899_395899 ; 
   reg __395899_395899;
   reg _395900_395900 ; 
   reg __395900_395900;
   reg _395901_395901 ; 
   reg __395901_395901;
   reg _395902_395902 ; 
   reg __395902_395902;
   reg _395903_395903 ; 
   reg __395903_395903;
   reg _395904_395904 ; 
   reg __395904_395904;
   reg _395905_395905 ; 
   reg __395905_395905;
   reg _395906_395906 ; 
   reg __395906_395906;
   reg _395907_395907 ; 
   reg __395907_395907;
   reg _395908_395908 ; 
   reg __395908_395908;
   reg _395909_395909 ; 
   reg __395909_395909;
   reg _395910_395910 ; 
   reg __395910_395910;
   reg _395911_395911 ; 
   reg __395911_395911;
   reg _395912_395912 ; 
   reg __395912_395912;
   reg _395913_395913 ; 
   reg __395913_395913;
   reg _395914_395914 ; 
   reg __395914_395914;
   reg _395915_395915 ; 
   reg __395915_395915;
   reg _395916_395916 ; 
   reg __395916_395916;
   reg _395917_395917 ; 
   reg __395917_395917;
   reg _395918_395918 ; 
   reg __395918_395918;
   reg _395919_395919 ; 
   reg __395919_395919;
   reg _395920_395920 ; 
   reg __395920_395920;
   reg _395921_395921 ; 
   reg __395921_395921;
   reg _395922_395922 ; 
   reg __395922_395922;
   reg _395923_395923 ; 
   reg __395923_395923;
   reg _395924_395924 ; 
   reg __395924_395924;
   reg _395925_395925 ; 
   reg __395925_395925;
   reg _395926_395926 ; 
   reg __395926_395926;
   reg _395927_395927 ; 
   reg __395927_395927;
   reg _395928_395928 ; 
   reg __395928_395928;
   reg _395929_395929 ; 
   reg __395929_395929;
   reg _395930_395930 ; 
   reg __395930_395930;
   reg _395931_395931 ; 
   reg __395931_395931;
   reg _395932_395932 ; 
   reg __395932_395932;
   reg _395933_395933 ; 
   reg __395933_395933;
   reg _395934_395934 ; 
   reg __395934_395934;
   reg _395935_395935 ; 
   reg __395935_395935;
   reg _395936_395936 ; 
   reg __395936_395936;
   reg _395937_395937 ; 
   reg __395937_395937;
   reg _395938_395938 ; 
   reg __395938_395938;
   reg _395939_395939 ; 
   reg __395939_395939;
   reg _395940_395940 ; 
   reg __395940_395940;
   reg _395941_395941 ; 
   reg __395941_395941;
   reg _395942_395942 ; 
   reg __395942_395942;
   reg _395943_395943 ; 
   reg __395943_395943;
   reg _395944_395944 ; 
   reg __395944_395944;
   reg _395945_395945 ; 
   reg __395945_395945;
   reg _395946_395946 ; 
   reg __395946_395946;
   reg _395947_395947 ; 
   reg __395947_395947;
   reg _395948_395948 ; 
   reg __395948_395948;
   reg _395949_395949 ; 
   reg __395949_395949;
   reg _395950_395950 ; 
   reg __395950_395950;
   reg _395951_395951 ; 
   reg __395951_395951;
   reg _395952_395952 ; 
   reg __395952_395952;
   reg _395953_395953 ; 
   reg __395953_395953;
   reg _395954_395954 ; 
   reg __395954_395954;
   reg _395955_395955 ; 
   reg __395955_395955;
   reg _395956_395956 ; 
   reg __395956_395956;
   reg _395957_395957 ; 
   reg __395957_395957;
   reg _395958_395958 ; 
   reg __395958_395958;
   reg _395959_395959 ; 
   reg __395959_395959;
   reg _395960_395960 ; 
   reg __395960_395960;
   reg _395961_395961 ; 
   reg __395961_395961;
   reg _395962_395962 ; 
   reg __395962_395962;
   reg _395963_395963 ; 
   reg __395963_395963;
   reg _395964_395964 ; 
   reg __395964_395964;
   reg _395965_395965 ; 
   reg __395965_395965;
   reg _395966_395966 ; 
   reg __395966_395966;
   reg _395967_395967 ; 
   reg __395967_395967;
   reg _395968_395968 ; 
   reg __395968_395968;
   reg _395969_395969 ; 
   reg __395969_395969;
   reg _395970_395970 ; 
   reg __395970_395970;
   reg _395971_395971 ; 
   reg __395971_395971;
   reg _395972_395972 ; 
   reg __395972_395972;
   reg _395973_395973 ; 
   reg __395973_395973;
   reg _395974_395974 ; 
   reg __395974_395974;
   reg _395975_395975 ; 
   reg __395975_395975;
   reg _395976_395976 ; 
   reg __395976_395976;
   reg _395977_395977 ; 
   reg __395977_395977;
   reg _395978_395978 ; 
   reg __395978_395978;
   reg _395979_395979 ; 
   reg __395979_395979;
   reg _395980_395980 ; 
   reg __395980_395980;
   reg _395981_395981 ; 
   reg __395981_395981;
   reg _395982_395982 ; 
   reg __395982_395982;
   reg _395983_395983 ; 
   reg __395983_395983;
   reg _395984_395984 ; 
   reg __395984_395984;
   reg _395985_395985 ; 
   reg __395985_395985;
   reg _395986_395986 ; 
   reg __395986_395986;
   reg _395987_395987 ; 
   reg __395987_395987;
   reg _395988_395988 ; 
   reg __395988_395988;
   reg _395989_395989 ; 
   reg __395989_395989;
   reg _395990_395990 ; 
   reg __395990_395990;
   reg _395991_395991 ; 
   reg __395991_395991;
   reg _395992_395992 ; 
   reg __395992_395992;
   reg _395993_395993 ; 
   reg __395993_395993;
   reg _395994_395994 ; 
   reg __395994_395994;
   reg _395995_395995 ; 
   reg __395995_395995;
   reg _395996_395996 ; 
   reg __395996_395996;
   reg _395997_395997 ; 
   reg __395997_395997;
   reg _395998_395998 ; 
   reg __395998_395998;
   reg _395999_395999 ; 
   reg __395999_395999;
   reg _396000_396000 ; 
   reg __396000_396000;
   reg _396001_396001 ; 
   reg __396001_396001;
   reg _396002_396002 ; 
   reg __396002_396002;
   reg _396003_396003 ; 
   reg __396003_396003;
   reg _396004_396004 ; 
   reg __396004_396004;
   reg _396005_396005 ; 
   reg __396005_396005;
   reg _396006_396006 ; 
   reg __396006_396006;
   reg _396007_396007 ; 
   reg __396007_396007;
   reg _396008_396008 ; 
   reg __396008_396008;
   reg _396009_396009 ; 
   reg __396009_396009;
   reg _396010_396010 ; 
   reg __396010_396010;
   reg _396011_396011 ; 
   reg __396011_396011;
   reg _396012_396012 ; 
   reg __396012_396012;
   reg _396013_396013 ; 
   reg __396013_396013;
   reg _396014_396014 ; 
   reg __396014_396014;
   reg _396015_396015 ; 
   reg __396015_396015;
   reg _396016_396016 ; 
   reg __396016_396016;
   reg _396017_396017 ; 
   reg __396017_396017;
   reg _396018_396018 ; 
   reg __396018_396018;
   reg _396019_396019 ; 
   reg __396019_396019;
   reg _396020_396020 ; 
   reg __396020_396020;
   reg _396021_396021 ; 
   reg __396021_396021;
   reg _396022_396022 ; 
   reg __396022_396022;
   reg _396023_396023 ; 
   reg __396023_396023;
   reg _396024_396024 ; 
   reg __396024_396024;
   reg _396025_396025 ; 
   reg __396025_396025;
   reg _396026_396026 ; 
   reg __396026_396026;
   reg _396027_396027 ; 
   reg __396027_396027;
   reg _396028_396028 ; 
   reg __396028_396028;
   reg _396029_396029 ; 
   reg __396029_396029;
   reg _396030_396030 ; 
   reg __396030_396030;
   reg _396031_396031 ; 
   reg __396031_396031;
   reg _396032_396032 ; 
   reg __396032_396032;
   reg _396033_396033 ; 
   reg __396033_396033;
   reg _396034_396034 ; 
   reg __396034_396034;
   reg _396035_396035 ; 
   reg __396035_396035;
   reg _396036_396036 ; 
   reg __396036_396036;
   reg _396037_396037 ; 
   reg __396037_396037;
   reg _396038_396038 ; 
   reg __396038_396038;
   reg _396039_396039 ; 
   reg __396039_396039;
   reg _396040_396040 ; 
   reg __396040_396040;
   reg _396041_396041 ; 
   reg __396041_396041;
   reg _396042_396042 ; 
   reg __396042_396042;
   reg _396043_396043 ; 
   reg __396043_396043;
   reg _396044_396044 ; 
   reg __396044_396044;
   reg _396045_396045 ; 
   reg __396045_396045;
   reg _396046_396046 ; 
   reg __396046_396046;
   reg _396047_396047 ; 
   reg __396047_396047;
   reg _396048_396048 ; 
   reg __396048_396048;
   reg _396049_396049 ; 
   reg __396049_396049;
   reg _396050_396050 ; 
   reg __396050_396050;
   reg _396051_396051 ; 
   reg __396051_396051;
   reg _396052_396052 ; 
   reg __396052_396052;
   reg _396053_396053 ; 
   reg __396053_396053;
   reg _396054_396054 ; 
   reg __396054_396054;
   reg _396055_396055 ; 
   reg __396055_396055;
   reg _396056_396056 ; 
   reg __396056_396056;
   reg _396057_396057 ; 
   reg __396057_396057;
   reg _396058_396058 ; 
   reg __396058_396058;
   reg _396059_396059 ; 
   reg __396059_396059;
   reg _396060_396060 ; 
   reg __396060_396060;
   reg _396061_396061 ; 
   reg __396061_396061;
   reg _396062_396062 ; 
   reg __396062_396062;
   reg _396063_396063 ; 
   reg __396063_396063;
   reg _396064_396064 ; 
   reg __396064_396064;
   reg _396065_396065 ; 
   reg __396065_396065;
   reg _396066_396066 ; 
   reg __396066_396066;
   reg _396067_396067 ; 
   reg __396067_396067;
   reg _396068_396068 ; 
   reg __396068_396068;
   reg _396069_396069 ; 
   reg __396069_396069;
   reg _396070_396070 ; 
   reg __396070_396070;
   reg _396071_396071 ; 
   reg __396071_396071;
   reg _396072_396072 ; 
   reg __396072_396072;
   reg _396073_396073 ; 
   reg __396073_396073;
   reg _396074_396074 ; 
   reg __396074_396074;
   reg _396075_396075 ; 
   reg __396075_396075;
   reg _396076_396076 ; 
   reg __396076_396076;
   reg _396077_396077 ; 
   reg __396077_396077;
   reg _396078_396078 ; 
   reg __396078_396078;
   reg _396079_396079 ; 
   reg __396079_396079;
   reg _396080_396080 ; 
   reg __396080_396080;
   reg _396081_396081 ; 
   reg __396081_396081;
   reg _396082_396082 ; 
   reg __396082_396082;
   reg _396083_396083 ; 
   reg __396083_396083;
   reg _396084_396084 ; 
   reg __396084_396084;
   reg _396085_396085 ; 
   reg __396085_396085;
   reg _396086_396086 ; 
   reg __396086_396086;
   reg _396087_396087 ; 
   reg __396087_396087;
   reg _396088_396088 ; 
   reg __396088_396088;
   reg _396089_396089 ; 
   reg __396089_396089;
   reg _396090_396090 ; 
   reg __396090_396090;
   reg _396091_396091 ; 
   reg __396091_396091;
   reg _396092_396092 ; 
   reg __396092_396092;
   reg _396093_396093 ; 
   reg __396093_396093;
   reg _396094_396094 ; 
   reg __396094_396094;
   reg _396095_396095 ; 
   reg __396095_396095;
   reg _396096_396096 ; 
   reg __396096_396096;
   reg _396097_396097 ; 
   reg __396097_396097;
   reg _396098_396098 ; 
   reg __396098_396098;
   reg _396099_396099 ; 
   reg __396099_396099;
   reg _396100_396100 ; 
   reg __396100_396100;
   reg _396101_396101 ; 
   reg __396101_396101;
   reg _396102_396102 ; 
   reg __396102_396102;
   reg _396103_396103 ; 
   reg __396103_396103;
   reg _396104_396104 ; 
   reg __396104_396104;
   reg _396105_396105 ; 
   reg __396105_396105;
   reg _396106_396106 ; 
   reg __396106_396106;
   reg _396107_396107 ; 
   reg __396107_396107;
   reg _396108_396108 ; 
   reg __396108_396108;
   reg _396109_396109 ; 
   reg __396109_396109;
   reg _396110_396110 ; 
   reg __396110_396110;
   reg _396111_396111 ; 
   reg __396111_396111;
   reg _396112_396112 ; 
   reg __396112_396112;
   reg _396113_396113 ; 
   reg __396113_396113;
   reg _396114_396114 ; 
   reg __396114_396114;
   reg _396115_396115 ; 
   reg __396115_396115;
   reg _396116_396116 ; 
   reg __396116_396116;
   reg _396117_396117 ; 
   reg __396117_396117;
   reg _396118_396118 ; 
   reg __396118_396118;
   reg _396119_396119 ; 
   reg __396119_396119;
   reg _396120_396120 ; 
   reg __396120_396120;
   reg _396121_396121 ; 
   reg __396121_396121;
   reg _396122_396122 ; 
   reg __396122_396122;
   reg _396123_396123 ; 
   reg __396123_396123;
   reg _396124_396124 ; 
   reg __396124_396124;
   reg _396125_396125 ; 
   reg __396125_396125;
   reg _396126_396126 ; 
   reg __396126_396126;
   reg _396127_396127 ; 
   reg __396127_396127;
   reg _396128_396128 ; 
   reg __396128_396128;
   reg _396129_396129 ; 
   reg __396129_396129;
   reg _396130_396130 ; 
   reg __396130_396130;
   reg _396131_396131 ; 
   reg __396131_396131;
   reg _396132_396132 ; 
   reg __396132_396132;
   reg _396133_396133 ; 
   reg __396133_396133;
   reg _396134_396134 ; 
   reg __396134_396134;
   reg _396135_396135 ; 
   reg __396135_396135;
   reg _396136_396136 ; 
   reg __396136_396136;
   reg _396137_396137 ; 
   reg __396137_396137;
   reg _396138_396138 ; 
   reg __396138_396138;
   reg _396139_396139 ; 
   reg __396139_396139;
   reg _396140_396140 ; 
   reg __396140_396140;
   reg _396141_396141 ; 
   reg __396141_396141;
   reg _396142_396142 ; 
   reg __396142_396142;
   reg _396143_396143 ; 
   reg __396143_396143;
   reg _396144_396144 ; 
   reg __396144_396144;
   reg _396145_396145 ; 
   reg __396145_396145;
   reg _396146_396146 ; 
   reg __396146_396146;
   reg _396147_396147 ; 
   reg __396147_396147;
   reg _396148_396148 ; 
   reg __396148_396148;
   reg _396149_396149 ; 
   reg __396149_396149;
   reg _396150_396150 ; 
   reg __396150_396150;
   reg _396151_396151 ; 
   reg __396151_396151;
   reg _396152_396152 ; 
   reg __396152_396152;
   reg _396153_396153 ; 
   reg __396153_396153;
   reg _396154_396154 ; 
   reg __396154_396154;
   reg _396155_396155 ; 
   reg __396155_396155;
   reg _396156_396156 ; 
   reg __396156_396156;
   reg _396157_396157 ; 
   reg __396157_396157;
   reg _396158_396158 ; 
   reg __396158_396158;
   reg _396159_396159 ; 
   reg __396159_396159;
   reg _396160_396160 ; 
   reg __396160_396160;
   reg _396161_396161 ; 
   reg __396161_396161;
   reg _396162_396162 ; 
   reg __396162_396162;
   reg _396163_396163 ; 
   reg __396163_396163;
   reg _396164_396164 ; 
   reg __396164_396164;
   reg _396165_396165 ; 
   reg __396165_396165;
   reg _396166_396166 ; 
   reg __396166_396166;
   reg _396167_396167 ; 
   reg __396167_396167;
   reg _396168_396168 ; 
   reg __396168_396168;
   reg _396169_396169 ; 
   reg __396169_396169;
   reg _396170_396170 ; 
   reg __396170_396170;
   reg _396171_396171 ; 
   reg __396171_396171;
   reg _396172_396172 ; 
   reg __396172_396172;
   reg _396173_396173 ; 
   reg __396173_396173;
   reg _396174_396174 ; 
   reg __396174_396174;
   reg _396175_396175 ; 
   reg __396175_396175;
   reg _396176_396176 ; 
   reg __396176_396176;
   reg _396177_396177 ; 
   reg __396177_396177;
   reg _396178_396178 ; 
   reg __396178_396178;
   reg _396179_396179 ; 
   reg __396179_396179;
   reg _396180_396180 ; 
   reg __396180_396180;
   reg _396181_396181 ; 
   reg __396181_396181;
   reg _396182_396182 ; 
   reg __396182_396182;
   reg _396183_396183 ; 
   reg __396183_396183;
   reg _396184_396184 ; 
   reg __396184_396184;
   reg _396185_396185 ; 
   reg __396185_396185;
   reg _396186_396186 ; 
   reg __396186_396186;
   reg _396187_396187 ; 
   reg __396187_396187;
   reg _396188_396188 ; 
   reg __396188_396188;
   reg _396189_396189 ; 
   reg __396189_396189;
   reg _396190_396190 ; 
   reg __396190_396190;
   reg _396191_396191 ; 
   reg __396191_396191;
   reg _396192_396192 ; 
   reg __396192_396192;
   reg _396193_396193 ; 
   reg __396193_396193;
   reg _396194_396194 ; 
   reg __396194_396194;
   reg _396195_396195 ; 
   reg __396195_396195;
   reg _396196_396196 ; 
   reg __396196_396196;
   reg _396197_396197 ; 
   reg __396197_396197;
   reg _396198_396198 ; 
   reg __396198_396198;
   reg _396199_396199 ; 
   reg __396199_396199;
   reg _396200_396200 ; 
   reg __396200_396200;
   reg _396201_396201 ; 
   reg __396201_396201;
   reg _396202_396202 ; 
   reg __396202_396202;
   reg _396203_396203 ; 
   reg __396203_396203;
   reg _396204_396204 ; 
   reg __396204_396204;
   reg _396205_396205 ; 
   reg __396205_396205;
   reg _396206_396206 ; 
   reg __396206_396206;
   reg _396207_396207 ; 
   reg __396207_396207;
   reg _396208_396208 ; 
   reg __396208_396208;
   reg _396209_396209 ; 
   reg __396209_396209;
   reg _396210_396210 ; 
   reg __396210_396210;
   reg _396211_396211 ; 
   reg __396211_396211;
   reg _396212_396212 ; 
   reg __396212_396212;
   reg _396213_396213 ; 
   reg __396213_396213;
   reg _396214_396214 ; 
   reg __396214_396214;
   reg _396215_396215 ; 
   reg __396215_396215;
   reg _396216_396216 ; 
   reg __396216_396216;
   reg _396217_396217 ; 
   reg __396217_396217;
   reg _396218_396218 ; 
   reg __396218_396218;
   reg _396219_396219 ; 
   reg __396219_396219;
   reg _396220_396220 ; 
   reg __396220_396220;
   reg _396221_396221 ; 
   reg __396221_396221;
   reg _396222_396222 ; 
   reg __396222_396222;
   reg _396223_396223 ; 
   reg __396223_396223;
   reg _396224_396224 ; 
   reg __396224_396224;
   reg _396225_396225 ; 
   reg __396225_396225;
   reg _396226_396226 ; 
   reg __396226_396226;
   reg _396227_396227 ; 
   reg __396227_396227;
   reg _396228_396228 ; 
   reg __396228_396228;
   reg _396229_396229 ; 
   reg __396229_396229;
   reg _396230_396230 ; 
   reg __396230_396230;
   reg _396231_396231 ; 
   reg __396231_396231;
   reg _396232_396232 ; 
   reg __396232_396232;
   reg _396233_396233 ; 
   reg __396233_396233;
   reg _396234_396234 ; 
   reg __396234_396234;
   reg _396235_396235 ; 
   reg __396235_396235;
   reg _396236_396236 ; 
   reg __396236_396236;
   reg _396237_396237 ; 
   reg __396237_396237;
   reg _396238_396238 ; 
   reg __396238_396238;
   reg _396239_396239 ; 
   reg __396239_396239;
   reg _396240_396240 ; 
   reg __396240_396240;
   reg _396241_396241 ; 
   reg __396241_396241;
   reg _396242_396242 ; 
   reg __396242_396242;
   reg _396243_396243 ; 
   reg __396243_396243;
   reg _396244_396244 ; 
   reg __396244_396244;
   reg _396245_396245 ; 
   reg __396245_396245;
   reg _396246_396246 ; 
   reg __396246_396246;
   reg _396247_396247 ; 
   reg __396247_396247;
   reg _396248_396248 ; 
   reg __396248_396248;
   reg _396249_396249 ; 
   reg __396249_396249;
   reg _396250_396250 ; 
   reg __396250_396250;
   reg _396251_396251 ; 
   reg __396251_396251;
   reg _396252_396252 ; 
   reg __396252_396252;
   reg _396253_396253 ; 
   reg __396253_396253;
   reg _396254_396254 ; 
   reg __396254_396254;
   reg _396255_396255 ; 
   reg __396255_396255;
   reg _396256_396256 ; 
   reg __396256_396256;
   reg _396257_396257 ; 
   reg __396257_396257;
   reg _396258_396258 ; 
   reg __396258_396258;
   reg _396259_396259 ; 
   reg __396259_396259;
   reg _396260_396260 ; 
   reg __396260_396260;
   reg _396261_396261 ; 
   reg __396261_396261;
   reg _396262_396262 ; 
   reg __396262_396262;
   reg _396263_396263 ; 
   reg __396263_396263;
   reg _396264_396264 ; 
   reg __396264_396264;
   reg _396265_396265 ; 
   reg __396265_396265;
   reg _396266_396266 ; 
   reg __396266_396266;
   reg _396267_396267 ; 
   reg __396267_396267;
   reg _396268_396268 ; 
   reg __396268_396268;
   reg _396269_396269 ; 
   reg __396269_396269;
   reg _396270_396270 ; 
   reg __396270_396270;
   reg _396271_396271 ; 
   reg __396271_396271;
   reg _396272_396272 ; 
   reg __396272_396272;
   reg _396273_396273 ; 
   reg __396273_396273;
   reg _396274_396274 ; 
   reg __396274_396274;
   reg _396275_396275 ; 
   reg __396275_396275;
   reg _396276_396276 ; 
   reg __396276_396276;
   reg _396277_396277 ; 
   reg __396277_396277;
   reg _396278_396278 ; 
   reg __396278_396278;
   reg _396279_396279 ; 
   reg __396279_396279;
   reg _396280_396280 ; 
   reg __396280_396280;
   reg _396281_396281 ; 
   reg __396281_396281;
   reg _396282_396282 ; 
   reg __396282_396282;
   reg _396283_396283 ; 
   reg __396283_396283;
   reg _396284_396284 ; 
   reg __396284_396284;
   reg _396285_396285 ; 
   reg __396285_396285;
   reg _396286_396286 ; 
   reg __396286_396286;
   reg _396287_396287 ; 
   reg __396287_396287;
   reg _396288_396288 ; 
   reg __396288_396288;
   reg _396289_396289 ; 
   reg __396289_396289;
   reg _396290_396290 ; 
   reg __396290_396290;
   reg _396291_396291 ; 
   reg __396291_396291;
   reg _396292_396292 ; 
   reg __396292_396292;
   reg _396293_396293 ; 
   reg __396293_396293;
   reg _396294_396294 ; 
   reg __396294_396294;
   reg _396295_396295 ; 
   reg __396295_396295;
   reg _396296_396296 ; 
   reg __396296_396296;
   reg _396297_396297 ; 
   reg __396297_396297;
   reg _396298_396298 ; 
   reg __396298_396298;
   reg _396299_396299 ; 
   reg __396299_396299;
   reg _396300_396300 ; 
   reg __396300_396300;
   reg _396301_396301 ; 
   reg __396301_396301;
   reg _396302_396302 ; 
   reg __396302_396302;
   reg _396303_396303 ; 
   reg __396303_396303;
   reg _396304_396304 ; 
   reg __396304_396304;
   reg _396305_396305 ; 
   reg __396305_396305;
   reg _396306_396306 ; 
   reg __396306_396306;
   reg _396307_396307 ; 
   reg __396307_396307;
   reg _396308_396308 ; 
   reg __396308_396308;
   reg _396309_396309 ; 
   reg __396309_396309;
   reg _396310_396310 ; 
   reg __396310_396310;
   reg _396311_396311 ; 
   reg __396311_396311;
   reg _396312_396312 ; 
   reg __396312_396312;
   reg _396313_396313 ; 
   reg __396313_396313;
   reg _396314_396314 ; 
   reg __396314_396314;
   reg _396315_396315 ; 
   reg __396315_396315;
   reg _396316_396316 ; 
   reg __396316_396316;
   reg _396317_396317 ; 
   reg __396317_396317;
   reg _396318_396318 ; 
   reg __396318_396318;
   reg _396319_396319 ; 
   reg __396319_396319;
   reg _396320_396320 ; 
   reg __396320_396320;
   reg _396321_396321 ; 
   reg __396321_396321;
   reg _396322_396322 ; 
   reg __396322_396322;
   reg _396323_396323 ; 
   reg __396323_396323;
   reg _396324_396324 ; 
   reg __396324_396324;
   reg _396325_396325 ; 
   reg __396325_396325;
   reg _396326_396326 ; 
   reg __396326_396326;
   reg _396327_396327 ; 
   reg __396327_396327;
   reg _396328_396328 ; 
   reg __396328_396328;
   reg _396329_396329 ; 
   reg __396329_396329;
   reg _396330_396330 ; 
   reg __396330_396330;
   reg _396331_396331 ; 
   reg __396331_396331;
   reg _396332_396332 ; 
   reg __396332_396332;
   reg _396333_396333 ; 
   reg __396333_396333;
   reg _396334_396334 ; 
   reg __396334_396334;
   reg _396335_396335 ; 
   reg __396335_396335;
   reg _396336_396336 ; 
   reg __396336_396336;
   reg _396337_396337 ; 
   reg __396337_396337;
   reg _396338_396338 ; 
   reg __396338_396338;
   reg _396339_396339 ; 
   reg __396339_396339;
   reg _396340_396340 ; 
   reg __396340_396340;
   reg _396341_396341 ; 
   reg __396341_396341;
   reg _396342_396342 ; 
   reg __396342_396342;
   reg _396343_396343 ; 
   reg __396343_396343;
   reg _396344_396344 ; 
   reg __396344_396344;
   reg _396345_396345 ; 
   reg __396345_396345;
   reg _396346_396346 ; 
   reg __396346_396346;
   reg _396347_396347 ; 
   reg __396347_396347;
   reg _396348_396348 ; 
   reg __396348_396348;
   reg _396349_396349 ; 
   reg __396349_396349;
   reg _396350_396350 ; 
   reg __396350_396350;
   reg _396351_396351 ; 
   reg __396351_396351;
   reg _396352_396352 ; 
   reg __396352_396352;
   reg _396353_396353 ; 
   reg __396353_396353;
   reg _396354_396354 ; 
   reg __396354_396354;
   reg _396355_396355 ; 
   reg __396355_396355;
   reg _396356_396356 ; 
   reg __396356_396356;
   reg _396357_396357 ; 
   reg __396357_396357;
   reg _396358_396358 ; 
   reg __396358_396358;
   reg _396359_396359 ; 
   reg __396359_396359;
   reg _396360_396360 ; 
   reg __396360_396360;
   reg _396361_396361 ; 
   reg __396361_396361;
   reg _396362_396362 ; 
   reg __396362_396362;
   reg _396363_396363 ; 
   reg __396363_396363;
   reg _396364_396364 ; 
   reg __396364_396364;
   reg _396365_396365 ; 
   reg __396365_396365;
   reg _396366_396366 ; 
   reg __396366_396366;
   reg _396367_396367 ; 
   reg __396367_396367;
   reg _396368_396368 ; 
   reg __396368_396368;
   reg _396369_396369 ; 
   reg __396369_396369;
   reg _396370_396370 ; 
   reg __396370_396370;
   reg _396371_396371 ; 
   reg __396371_396371;
   reg _396372_396372 ; 
   reg __396372_396372;
   reg _396373_396373 ; 
   reg __396373_396373;
   reg _396374_396374 ; 
   reg __396374_396374;
   reg _396375_396375 ; 
   reg __396375_396375;
   reg _396376_396376 ; 
   reg __396376_396376;
   reg _396377_396377 ; 
   reg __396377_396377;
   reg _396378_396378 ; 
   reg __396378_396378;
   reg _396379_396379 ; 
   reg __396379_396379;
   reg _396380_396380 ; 
   reg __396380_396380;
   reg _396381_396381 ; 
   reg __396381_396381;
   reg _396382_396382 ; 
   reg __396382_396382;
   reg _396383_396383 ; 
   reg __396383_396383;
   reg _396384_396384 ; 
   reg __396384_396384;
   reg _396385_396385 ; 
   reg __396385_396385;
   reg _396386_396386 ; 
   reg __396386_396386;
   reg _396387_396387 ; 
   reg __396387_396387;
   reg _396388_396388 ; 
   reg __396388_396388;
   reg _396389_396389 ; 
   reg __396389_396389;
   reg _396390_396390 ; 
   reg __396390_396390;
   reg _396391_396391 ; 
   reg __396391_396391;
   reg _396392_396392 ; 
   reg __396392_396392;
   reg _396393_396393 ; 
   reg __396393_396393;
   reg _396394_396394 ; 
   reg __396394_396394;
   reg _396395_396395 ; 
   reg __396395_396395;
   reg _396396_396396 ; 
   reg __396396_396396;
   reg _396397_396397 ; 
   reg __396397_396397;
   reg _396398_396398 ; 
   reg __396398_396398;
   reg _396399_396399 ; 
   reg __396399_396399;
   reg _396400_396400 ; 
   reg __396400_396400;
   reg _396401_396401 ; 
   reg __396401_396401;
   reg _396402_396402 ; 
   reg __396402_396402;
   reg _396403_396403 ; 
   reg __396403_396403;
   reg _396404_396404 ; 
   reg __396404_396404;
   reg _396405_396405 ; 
   reg __396405_396405;
   reg _396406_396406 ; 
   reg __396406_396406;
   reg _396407_396407 ; 
   reg __396407_396407;
   reg _396408_396408 ; 
   reg __396408_396408;
   reg _396409_396409 ; 
   reg __396409_396409;
   reg _396410_396410 ; 
   reg __396410_396410;
   reg _396411_396411 ; 
   reg __396411_396411;
   reg _396412_396412 ; 
   reg __396412_396412;
   reg _396413_396413 ; 
   reg __396413_396413;
   reg _396414_396414 ; 
   reg __396414_396414;
   reg _396415_396415 ; 
   reg __396415_396415;
   reg _396416_396416 ; 
   reg __396416_396416;
   reg _396417_396417 ; 
   reg __396417_396417;
   reg _396418_396418 ; 
   reg __396418_396418;
   reg _396419_396419 ; 
   reg __396419_396419;
   reg _396420_396420 ; 
   reg __396420_396420;
   reg _396421_396421 ; 
   reg __396421_396421;
   reg _396422_396422 ; 
   reg __396422_396422;
   reg _396423_396423 ; 
   reg __396423_396423;
   reg _396424_396424 ; 
   reg __396424_396424;
   reg _396425_396425 ; 
   reg __396425_396425;
   reg _396426_396426 ; 
   reg __396426_396426;
   reg _396427_396427 ; 
   reg __396427_396427;
   reg _396428_396428 ; 
   reg __396428_396428;
   reg _396429_396429 ; 
   reg __396429_396429;
   reg _396430_396430 ; 
   reg __396430_396430;
   reg _396431_396431 ; 
   reg __396431_396431;
   reg _396432_396432 ; 
   reg __396432_396432;
   reg _396433_396433 ; 
   reg __396433_396433;
   reg _396434_396434 ; 
   reg __396434_396434;
   reg _396435_396435 ; 
   reg __396435_396435;
   reg _396436_396436 ; 
   reg __396436_396436;
   reg _396437_396437 ; 
   reg __396437_396437;
   reg _396438_396438 ; 
   reg __396438_396438;
   reg _396439_396439 ; 
   reg __396439_396439;
   reg _396440_396440 ; 
   reg __396440_396440;
   reg _396441_396441 ; 
   reg __396441_396441;
   reg _396442_396442 ; 
   reg __396442_396442;
   reg _396443_396443 ; 
   reg __396443_396443;
   reg _396444_396444 ; 
   reg __396444_396444;
   reg _396445_396445 ; 
   reg __396445_396445;
   reg _396446_396446 ; 
   reg __396446_396446;
   reg _396447_396447 ; 
   reg __396447_396447;
   reg _396448_396448 ; 
   reg __396448_396448;
   reg _396449_396449 ; 
   reg __396449_396449;
   reg _396450_396450 ; 
   reg __396450_396450;
   reg _396451_396451 ; 
   reg __396451_396451;
   reg _396452_396452 ; 
   reg __396452_396452;
   reg _396453_396453 ; 
   reg __396453_396453;
   reg _396454_396454 ; 
   reg __396454_396454;
   reg _396455_396455 ; 
   reg __396455_396455;
   reg _396456_396456 ; 
   reg __396456_396456;
   reg _396457_396457 ; 
   reg __396457_396457;
   reg _396458_396458 ; 
   reg __396458_396458;
   reg _396459_396459 ; 
   reg __396459_396459;
   reg _396460_396460 ; 
   reg __396460_396460;
   reg _396461_396461 ; 
   reg __396461_396461;
   reg _396462_396462 ; 
   reg __396462_396462;
   reg _396463_396463 ; 
   reg __396463_396463;
   reg _396464_396464 ; 
   reg __396464_396464;
   reg _396465_396465 ; 
   reg __396465_396465;
   reg _396466_396466 ; 
   reg __396466_396466;
   reg _396467_396467 ; 
   reg __396467_396467;
   reg _396468_396468 ; 
   reg __396468_396468;
   reg _396469_396469 ; 
   reg __396469_396469;
   reg _396470_396470 ; 
   reg __396470_396470;
   reg _396471_396471 ; 
   reg __396471_396471;
   reg _396472_396472 ; 
   reg __396472_396472;
   reg _396473_396473 ; 
   reg __396473_396473;
   reg _396474_396474 ; 
   reg __396474_396474;
   reg _396475_396475 ; 
   reg __396475_396475;
   reg _396476_396476 ; 
   reg __396476_396476;
   reg _396477_396477 ; 
   reg __396477_396477;
   reg _396478_396478 ; 
   reg __396478_396478;
   reg _396479_396479 ; 
   reg __396479_396479;
   reg _396480_396480 ; 
   reg __396480_396480;
   reg _396481_396481 ; 
   reg __396481_396481;
   reg _396482_396482 ; 
   reg __396482_396482;
   reg _396483_396483 ; 
   reg __396483_396483;
   reg _396484_396484 ; 
   reg __396484_396484;
   reg _396485_396485 ; 
   reg __396485_396485;
   reg _396486_396486 ; 
   reg __396486_396486;
   reg _396487_396487 ; 
   reg __396487_396487;
   reg _396488_396488 ; 
   reg __396488_396488;
   reg _396489_396489 ; 
   reg __396489_396489;
   reg _396490_396490 ; 
   reg __396490_396490;
   reg _396491_396491 ; 
   reg __396491_396491;
   reg _396492_396492 ; 
   reg __396492_396492;
   reg _396493_396493 ; 
   reg __396493_396493;
   reg _396494_396494 ; 
   reg __396494_396494;
   reg _396495_396495 ; 
   reg __396495_396495;
   reg _396496_396496 ; 
   reg __396496_396496;
   reg _396497_396497 ; 
   reg __396497_396497;
   reg _396498_396498 ; 
   reg __396498_396498;
   reg _396499_396499 ; 
   reg __396499_396499;
   reg _396500_396500 ; 
   reg __396500_396500;
   reg _396501_396501 ; 
   reg __396501_396501;
   reg _396502_396502 ; 
   reg __396502_396502;
   reg _396503_396503 ; 
   reg __396503_396503;
   reg _396504_396504 ; 
   reg __396504_396504;
   reg _396505_396505 ; 
   reg __396505_396505;
   reg _396506_396506 ; 
   reg __396506_396506;
   reg _396507_396507 ; 
   reg __396507_396507;
   reg _396508_396508 ; 
   reg __396508_396508;
   reg _396509_396509 ; 
   reg __396509_396509;
   reg _396510_396510 ; 
   reg __396510_396510;
   reg _396511_396511 ; 
   reg __396511_396511;
   reg _396512_396512 ; 
   reg __396512_396512;
   reg _396513_396513 ; 
   reg __396513_396513;
   reg _396514_396514 ; 
   reg __396514_396514;
   reg _396515_396515 ; 
   reg __396515_396515;
   reg _396516_396516 ; 
   reg __396516_396516;
   reg _396517_396517 ; 
   reg __396517_396517;
   reg _396518_396518 ; 
   reg __396518_396518;
   reg _396519_396519 ; 
   reg __396519_396519;
   reg _396520_396520 ; 
   reg __396520_396520;
   reg _396521_396521 ; 
   reg __396521_396521;
   reg _396522_396522 ; 
   reg __396522_396522;
   reg _396523_396523 ; 
   reg __396523_396523;
   reg _396524_396524 ; 
   reg __396524_396524;
   reg _396525_396525 ; 
   reg __396525_396525;
   reg _396526_396526 ; 
   reg __396526_396526;
   reg _396527_396527 ; 
   reg __396527_396527;
   reg _396528_396528 ; 
   reg __396528_396528;
   reg _396529_396529 ; 
   reg __396529_396529;
   reg _396530_396530 ; 
   reg __396530_396530;
   reg _396531_396531 ; 
   reg __396531_396531;
   reg _396532_396532 ; 
   reg __396532_396532;
   reg _396533_396533 ; 
   reg __396533_396533;
   reg _396534_396534 ; 
   reg __396534_396534;
   reg _396535_396535 ; 
   reg __396535_396535;
   reg _396536_396536 ; 
   reg __396536_396536;
   reg _396537_396537 ; 
   reg __396537_396537;
   reg _396538_396538 ; 
   reg __396538_396538;
   reg _396539_396539 ; 
   reg __396539_396539;
   reg _396540_396540 ; 
   reg __396540_396540;
   reg _396541_396541 ; 
   reg __396541_396541;
   reg _396542_396542 ; 
   reg __396542_396542;
   reg _396543_396543 ; 
   reg __396543_396543;
   reg _396544_396544 ; 
   reg __396544_396544;
   reg _396545_396545 ; 
   reg __396545_396545;
   reg _396546_396546 ; 
   reg __396546_396546;
   reg _396547_396547 ; 
   reg __396547_396547;
   reg _396548_396548 ; 
   reg __396548_396548;
   reg _396549_396549 ; 
   reg __396549_396549;
   reg _396550_396550 ; 
   reg __396550_396550;
   reg _396551_396551 ; 
   reg __396551_396551;
   reg _396552_396552 ; 
   reg __396552_396552;
   reg _396553_396553 ; 
   reg __396553_396553;
   reg _396554_396554 ; 
   reg __396554_396554;
   reg _396555_396555 ; 
   reg __396555_396555;
   reg _396556_396556 ; 
   reg __396556_396556;
   reg _396557_396557 ; 
   reg __396557_396557;
   reg _396558_396558 ; 
   reg __396558_396558;
   reg _396559_396559 ; 
   reg __396559_396559;
   reg _396560_396560 ; 
   reg __396560_396560;
   reg _396561_396561 ; 
   reg __396561_396561;
   reg _396562_396562 ; 
   reg __396562_396562;
   reg _396563_396563 ; 
   reg __396563_396563;
   reg _396564_396564 ; 
   reg __396564_396564;
   reg _396565_396565 ; 
   reg __396565_396565;
   reg _396566_396566 ; 
   reg __396566_396566;
   reg _396567_396567 ; 
   reg __396567_396567;
   reg _396568_396568 ; 
   reg __396568_396568;
   reg _396569_396569 ; 
   reg __396569_396569;
   reg _396570_396570 ; 
   reg __396570_396570;
   reg _396571_396571 ; 
   reg __396571_396571;
   reg _396572_396572 ; 
   reg __396572_396572;
   reg _396573_396573 ; 
   reg __396573_396573;
   reg _396574_396574 ; 
   reg __396574_396574;
   reg _396575_396575 ; 
   reg __396575_396575;
   reg _396576_396576 ; 
   reg __396576_396576;
   reg _396577_396577 ; 
   reg __396577_396577;
   reg _396578_396578 ; 
   reg __396578_396578;
   reg _396579_396579 ; 
   reg __396579_396579;
   reg _396580_396580 ; 
   reg __396580_396580;
   reg _396581_396581 ; 
   reg __396581_396581;
   reg _396582_396582 ; 
   reg __396582_396582;
   reg _396583_396583 ; 
   reg __396583_396583;
   reg _396584_396584 ; 
   reg __396584_396584;
   reg _396585_396585 ; 
   reg __396585_396585;
   reg _396586_396586 ; 
   reg __396586_396586;
   reg _396587_396587 ; 
   reg __396587_396587;
   reg _396588_396588 ; 
   reg __396588_396588;
   reg _396589_396589 ; 
   reg __396589_396589;
   reg _396590_396590 ; 
   reg __396590_396590;
   reg _396591_396591 ; 
   reg __396591_396591;
   reg _396592_396592 ; 
   reg __396592_396592;
   reg _396593_396593 ; 
   reg __396593_396593;
   reg _396594_396594 ; 
   reg __396594_396594;
   reg _396595_396595 ; 
   reg __396595_396595;
   reg _396596_396596 ; 
   reg __396596_396596;
   reg _396597_396597 ; 
   reg __396597_396597;
   reg _396598_396598 ; 
   reg __396598_396598;
   reg _396599_396599 ; 
   reg __396599_396599;
   reg _396600_396600 ; 
   reg __396600_396600;
   reg _396601_396601 ; 
   reg __396601_396601;
   reg _396602_396602 ; 
   reg __396602_396602;
   reg _396603_396603 ; 
   reg __396603_396603;
   reg _396604_396604 ; 
   reg __396604_396604;
   reg _396605_396605 ; 
   reg __396605_396605;
   reg _396606_396606 ; 
   reg __396606_396606;
   reg _396607_396607 ; 
   reg __396607_396607;
   reg _396608_396608 ; 
   reg __396608_396608;
   reg _396609_396609 ; 
   reg __396609_396609;
   reg _396610_396610 ; 
   reg __396610_396610;
   reg _396611_396611 ; 
   reg __396611_396611;
   reg _396612_396612 ; 
   reg __396612_396612;
   reg _396613_396613 ; 
   reg __396613_396613;
   reg _396614_396614 ; 
   reg __396614_396614;
   reg _396615_396615 ; 
   reg __396615_396615;
   reg _396616_396616 ; 
   reg __396616_396616;
   reg _396617_396617 ; 
   reg __396617_396617;
   reg _396618_396618 ; 
   reg __396618_396618;
   reg _396619_396619 ; 
   reg __396619_396619;
   reg _396620_396620 ; 
   reg __396620_396620;
   reg _396621_396621 ; 
   reg __396621_396621;
   reg _396622_396622 ; 
   reg __396622_396622;
   reg _396623_396623 ; 
   reg __396623_396623;
   reg _396624_396624 ; 
   reg __396624_396624;
   reg _396625_396625 ; 
   reg __396625_396625;
   reg _396626_396626 ; 
   reg __396626_396626;
   reg _396627_396627 ; 
   reg __396627_396627;
   reg _396628_396628 ; 
   reg __396628_396628;
   reg _396629_396629 ; 
   reg __396629_396629;
   reg _396630_396630 ; 
   reg __396630_396630;
   reg _396631_396631 ; 
   reg __396631_396631;
   reg _396632_396632 ; 
   reg __396632_396632;
   reg _396633_396633 ; 
   reg __396633_396633;
   reg _396634_396634 ; 
   reg __396634_396634;
   reg _396635_396635 ; 
   reg __396635_396635;
   reg _396636_396636 ; 
   reg __396636_396636;
   reg _396637_396637 ; 
   reg __396637_396637;
   reg _396638_396638 ; 
   reg __396638_396638;
   reg _396639_396639 ; 
   reg __396639_396639;
   reg _396640_396640 ; 
   reg __396640_396640;
   reg _396641_396641 ; 
   reg __396641_396641;
   reg _396642_396642 ; 
   reg __396642_396642;
   reg _396643_396643 ; 
   reg __396643_396643;
   reg _396644_396644 ; 
   reg __396644_396644;
   reg _396645_396645 ; 
   reg __396645_396645;
   reg _396646_396646 ; 
   reg __396646_396646;
   reg _396647_396647 ; 
   reg __396647_396647;
   reg _396648_396648 ; 
   reg __396648_396648;
   reg _396649_396649 ; 
   reg __396649_396649;
   reg _396650_396650 ; 
   reg __396650_396650;
   reg _396651_396651 ; 
   reg __396651_396651;
   reg _396652_396652 ; 
   reg __396652_396652;
   reg _396653_396653 ; 
   reg __396653_396653;
   reg _396654_396654 ; 
   reg __396654_396654;
   reg _396655_396655 ; 
   reg __396655_396655;
   reg _396656_396656 ; 
   reg __396656_396656;
   reg _396657_396657 ; 
   reg __396657_396657;
   reg _396658_396658 ; 
   reg __396658_396658;
   reg _396659_396659 ; 
   reg __396659_396659;
   reg _396660_396660 ; 
   reg __396660_396660;
   reg _396661_396661 ; 
   reg __396661_396661;
   reg _396662_396662 ; 
   reg __396662_396662;
   reg _396663_396663 ; 
   reg __396663_396663;
   reg _396664_396664 ; 
   reg __396664_396664;
   reg _396665_396665 ; 
   reg __396665_396665;
   reg _396666_396666 ; 
   reg __396666_396666;
   reg _396667_396667 ; 
   reg __396667_396667;
   reg _396668_396668 ; 
   reg __396668_396668;
   reg _396669_396669 ; 
   reg __396669_396669;
   reg _396670_396670 ; 
   reg __396670_396670;
   reg _396671_396671 ; 
   reg __396671_396671;
   reg _396672_396672 ; 
   reg __396672_396672;
   reg _396673_396673 ; 
   reg __396673_396673;
   reg _396674_396674 ; 
   reg __396674_396674;
   reg _396675_396675 ; 
   reg __396675_396675;
   reg _396676_396676 ; 
   reg __396676_396676;
   reg _396677_396677 ; 
   reg __396677_396677;
   reg _396678_396678 ; 
   reg __396678_396678;
   reg _396679_396679 ; 
   reg __396679_396679;
   reg _396680_396680 ; 
   reg __396680_396680;
   reg _396681_396681 ; 
   reg __396681_396681;
   reg _396682_396682 ; 
   reg __396682_396682;
   reg _396683_396683 ; 
   reg __396683_396683;
   reg _396684_396684 ; 
   reg __396684_396684;
   reg _396685_396685 ; 
   reg __396685_396685;
   reg _396686_396686 ; 
   reg __396686_396686;
   reg _396687_396687 ; 
   reg __396687_396687;
   reg _396688_396688 ; 
   reg __396688_396688;
   reg _396689_396689 ; 
   reg __396689_396689;
   reg _396690_396690 ; 
   reg __396690_396690;
   reg _396691_396691 ; 
   reg __396691_396691;
   reg _396692_396692 ; 
   reg __396692_396692;
   reg _396693_396693 ; 
   reg __396693_396693;
   reg _396694_396694 ; 
   reg __396694_396694;
   reg _396695_396695 ; 
   reg __396695_396695;
   reg _396696_396696 ; 
   reg __396696_396696;
   reg _396697_396697 ; 
   reg __396697_396697;
   reg _396698_396698 ; 
   reg __396698_396698;
   reg _396699_396699 ; 
   reg __396699_396699;
   reg _396700_396700 ; 
   reg __396700_396700;
   reg _396701_396701 ; 
   reg __396701_396701;
   reg _396702_396702 ; 
   reg __396702_396702;
   reg _396703_396703 ; 
   reg __396703_396703;
   reg _396704_396704 ; 
   reg __396704_396704;
   reg _396705_396705 ; 
   reg __396705_396705;
   reg _396706_396706 ; 
   reg __396706_396706;
   reg _396707_396707 ; 
   reg __396707_396707;
   reg _396708_396708 ; 
   reg __396708_396708;
   reg _396709_396709 ; 
   reg __396709_396709;
   reg _396710_396710 ; 
   reg __396710_396710;
   reg _396711_396711 ; 
   reg __396711_396711;
   reg _396712_396712 ; 
   reg __396712_396712;
   reg _396713_396713 ; 
   reg __396713_396713;
   reg _396714_396714 ; 
   reg __396714_396714;
   reg _396715_396715 ; 
   reg __396715_396715;
   reg _396716_396716 ; 
   reg __396716_396716;
   reg _396717_396717 ; 
   reg __396717_396717;
   reg _396718_396718 ; 
   reg __396718_396718;
   reg _396719_396719 ; 
   reg __396719_396719;
   reg _396720_396720 ; 
   reg __396720_396720;
   reg _396721_396721 ; 
   reg __396721_396721;
   reg _396722_396722 ; 
   reg __396722_396722;
   reg _396723_396723 ; 
   reg __396723_396723;
   reg _396724_396724 ; 
   reg __396724_396724;
   reg _396725_396725 ; 
   reg __396725_396725;
   reg _396726_396726 ; 
   reg __396726_396726;
   reg _396727_396727 ; 
   reg __396727_396727;
   reg _396728_396728 ; 
   reg __396728_396728;
   reg _396729_396729 ; 
   reg __396729_396729;
   reg _396730_396730 ; 
   reg __396730_396730;
   reg _396731_396731 ; 
   reg __396731_396731;
   reg _396732_396732 ; 
   reg __396732_396732;
   reg _396733_396733 ; 
   reg __396733_396733;
   reg _396734_396734 ; 
   reg __396734_396734;
   reg _396735_396735 ; 
   reg __396735_396735;
   reg _396736_396736 ; 
   reg __396736_396736;
   reg _396737_396737 ; 
   reg __396737_396737;
   reg _396738_396738 ; 
   reg __396738_396738;
   reg _396739_396739 ; 
   reg __396739_396739;
   reg _396740_396740 ; 
   reg __396740_396740;
   reg _396741_396741 ; 
   reg __396741_396741;
   reg _396742_396742 ; 
   reg __396742_396742;
   reg _396743_396743 ; 
   reg __396743_396743;
   reg _396744_396744 ; 
   reg __396744_396744;
   reg _396745_396745 ; 
   reg __396745_396745;
   reg _396746_396746 ; 
   reg __396746_396746;
   reg _396747_396747 ; 
   reg __396747_396747;
   reg _396748_396748 ; 
   reg __396748_396748;
   reg _396749_396749 ; 
   reg __396749_396749;
   reg _396750_396750 ; 
   reg __396750_396750;
   reg _396751_396751 ; 
   reg __396751_396751;
   reg _396752_396752 ; 
   reg __396752_396752;
   reg _396753_396753 ; 
   reg __396753_396753;
   reg _396754_396754 ; 
   reg __396754_396754;
   reg _396755_396755 ; 
   reg __396755_396755;
   reg _396756_396756 ; 
   reg __396756_396756;
   reg _396757_396757 ; 
   reg __396757_396757;
   reg _396758_396758 ; 
   reg __396758_396758;
   reg _396759_396759 ; 
   reg __396759_396759;
   reg _396760_396760 ; 
   reg __396760_396760;
   reg _396761_396761 ; 
   reg __396761_396761;
   reg _396762_396762 ; 
   reg __396762_396762;
   reg _396763_396763 ; 
   reg __396763_396763;
   reg _396764_396764 ; 
   reg __396764_396764;
   reg _396765_396765 ; 
   reg __396765_396765;
   reg _396766_396766 ; 
   reg __396766_396766;
   reg _396767_396767 ; 
   reg __396767_396767;
   reg _396768_396768 ; 
   reg __396768_396768;
   reg _396769_396769 ; 
   reg __396769_396769;
   reg _396770_396770 ; 
   reg __396770_396770;
   reg _396771_396771 ; 
   reg __396771_396771;
   reg _396772_396772 ; 
   reg __396772_396772;
   reg _396773_396773 ; 
   reg __396773_396773;
   reg _396774_396774 ; 
   reg __396774_396774;
   reg _396775_396775 ; 
   reg __396775_396775;
   reg _396776_396776 ; 
   reg __396776_396776;
   reg _396777_396777 ; 
   reg __396777_396777;
   reg _396778_396778 ; 
   reg __396778_396778;
   reg _396779_396779 ; 
   reg __396779_396779;
   reg _396780_396780 ; 
   reg __396780_396780;
   reg _396781_396781 ; 
   reg __396781_396781;
   reg _396782_396782 ; 
   reg __396782_396782;
   reg _396783_396783 ; 
   reg __396783_396783;
   reg _396784_396784 ; 
   reg __396784_396784;
   reg _396785_396785 ; 
   reg __396785_396785;
   reg _396786_396786 ; 
   reg __396786_396786;
   reg _396787_396787 ; 
   reg __396787_396787;
   reg _396788_396788 ; 
   reg __396788_396788;
   reg _396789_396789 ; 
   reg __396789_396789;
   reg _396790_396790 ; 
   reg __396790_396790;
   reg _396791_396791 ; 
   reg __396791_396791;
   reg _396792_396792 ; 
   reg __396792_396792;
   reg _396793_396793 ; 
   reg __396793_396793;
   reg _396794_396794 ; 
   reg __396794_396794;
   reg _396795_396795 ; 
   reg __396795_396795;
   reg _396796_396796 ; 
   reg __396796_396796;
   reg _396797_396797 ; 
   reg __396797_396797;
   reg _396798_396798 ; 
   reg __396798_396798;
   reg _396799_396799 ; 
   reg __396799_396799;
   reg _396800_396800 ; 
   reg __396800_396800;
   reg _396801_396801 ; 
   reg __396801_396801;
   reg _396802_396802 ; 
   reg __396802_396802;
   reg _396803_396803 ; 
   reg __396803_396803;
   reg _396804_396804 ; 
   reg __396804_396804;
   reg _396805_396805 ; 
   reg __396805_396805;
   reg _396806_396806 ; 
   reg __396806_396806;
   reg _396807_396807 ; 
   reg __396807_396807;
   reg _396808_396808 ; 
   reg __396808_396808;
   reg _396809_396809 ; 
   reg __396809_396809;
   reg _396810_396810 ; 
   reg __396810_396810;
   reg _396811_396811 ; 
   reg __396811_396811;
   reg _396812_396812 ; 
   reg __396812_396812;
   reg _396813_396813 ; 
   reg __396813_396813;
   reg _396814_396814 ; 
   reg __396814_396814;
   reg _396815_396815 ; 
   reg __396815_396815;
   reg _396816_396816 ; 
   reg __396816_396816;
   reg _396817_396817 ; 
   reg __396817_396817;
   reg _396818_396818 ; 
   reg __396818_396818;
   reg _396819_396819 ; 
   reg __396819_396819;
   reg _396820_396820 ; 
   reg __396820_396820;
   reg _396821_396821 ; 
   reg __396821_396821;
   reg _396822_396822 ; 
   reg __396822_396822;
   reg _396823_396823 ; 
   reg __396823_396823;
   reg _396824_396824 ; 
   reg __396824_396824;
   reg _396825_396825 ; 
   reg __396825_396825;
   reg _396826_396826 ; 
   reg __396826_396826;
   reg _396827_396827 ; 
   reg __396827_396827;
   reg _396828_396828 ; 
   reg __396828_396828;
   reg _396829_396829 ; 
   reg __396829_396829;
   reg _396830_396830 ; 
   reg __396830_396830;
   reg _396831_396831 ; 
   reg __396831_396831;
   reg _396832_396832 ; 
   reg __396832_396832;
   reg _396833_396833 ; 
   reg __396833_396833;
   reg _396834_396834 ; 
   reg __396834_396834;
   reg _396835_396835 ; 
   reg __396835_396835;
   reg _396836_396836 ; 
   reg __396836_396836;
   reg _396837_396837 ; 
   reg __396837_396837;
   reg _396838_396838 ; 
   reg __396838_396838;
   reg _396839_396839 ; 
   reg __396839_396839;
   reg _396840_396840 ; 
   reg __396840_396840;
   reg _396841_396841 ; 
   reg __396841_396841;
   reg _396842_396842 ; 
   reg __396842_396842;
   reg _396843_396843 ; 
   reg __396843_396843;
   reg _396844_396844 ; 
   reg __396844_396844;
   reg _396845_396845 ; 
   reg __396845_396845;
   reg _396846_396846 ; 
   reg __396846_396846;
   reg _396847_396847 ; 
   reg __396847_396847;
   reg _396848_396848 ; 
   reg __396848_396848;
   reg _396849_396849 ; 
   reg __396849_396849;
   reg _396850_396850 ; 
   reg __396850_396850;
   reg _396851_396851 ; 
   reg __396851_396851;
   reg _396852_396852 ; 
   reg __396852_396852;
   reg _396853_396853 ; 
   reg __396853_396853;
   reg _396854_396854 ; 
   reg __396854_396854;
   reg _396855_396855 ; 
   reg __396855_396855;
   reg _396856_396856 ; 
   reg __396856_396856;
   reg _396857_396857 ; 
   reg __396857_396857;
   reg _396858_396858 ; 
   reg __396858_396858;
   reg _396859_396859 ; 
   reg __396859_396859;
   reg _396860_396860 ; 
   reg __396860_396860;
   reg _396861_396861 ; 
   reg __396861_396861;
   reg _396862_396862 ; 
   reg __396862_396862;
   reg _396863_396863 ; 
   reg __396863_396863;
   reg _396864_396864 ; 
   reg __396864_396864;
   reg _396865_396865 ; 
   reg __396865_396865;
   reg _396866_396866 ; 
   reg __396866_396866;
   reg _396867_396867 ; 
   reg __396867_396867;
   reg _396868_396868 ; 
   reg __396868_396868;
   reg _396869_396869 ; 
   reg __396869_396869;
   reg _396870_396870 ; 
   reg __396870_396870;
   reg _396871_396871 ; 
   reg __396871_396871;
   reg _396872_396872 ; 
   reg __396872_396872;
   reg _396873_396873 ; 
   reg __396873_396873;
   reg _396874_396874 ; 
   reg __396874_396874;
   reg _396875_396875 ; 
   reg __396875_396875;
   reg _396876_396876 ; 
   reg __396876_396876;
   reg _396877_396877 ; 
   reg __396877_396877;
   reg _396878_396878 ; 
   reg __396878_396878;
   reg _396879_396879 ; 
   reg __396879_396879;
   reg _396880_396880 ; 
   reg __396880_396880;
   reg _396881_396881 ; 
   reg __396881_396881;
   reg _396882_396882 ; 
   reg __396882_396882;
   reg _396883_396883 ; 
   reg __396883_396883;
   reg _396884_396884 ; 
   reg __396884_396884;
   reg _396885_396885 ; 
   reg __396885_396885;
   reg _396886_396886 ; 
   reg __396886_396886;
   reg _396887_396887 ; 
   reg __396887_396887;
   reg _396888_396888 ; 
   reg __396888_396888;
   reg _396889_396889 ; 
   reg __396889_396889;
   reg _396890_396890 ; 
   reg __396890_396890;
   reg _396891_396891 ; 
   reg __396891_396891;
   reg _396892_396892 ; 
   reg __396892_396892;
   reg _396893_396893 ; 
   reg __396893_396893;
   reg _396894_396894 ; 
   reg __396894_396894;
   reg _396895_396895 ; 
   reg __396895_396895;
   reg _396896_396896 ; 
   reg __396896_396896;
   reg _396897_396897 ; 
   reg __396897_396897;
   reg _396898_396898 ; 
   reg __396898_396898;
   reg _396899_396899 ; 
   reg __396899_396899;
   reg _396900_396900 ; 
   reg __396900_396900;
   reg _396901_396901 ; 
   reg __396901_396901;
   reg _396902_396902 ; 
   reg __396902_396902;
   reg _396903_396903 ; 
   reg __396903_396903;
   reg _396904_396904 ; 
   reg __396904_396904;
   reg _396905_396905 ; 
   reg __396905_396905;
   reg _396906_396906 ; 
   reg __396906_396906;
   reg _396907_396907 ; 
   reg __396907_396907;
   reg _396908_396908 ; 
   reg __396908_396908;
   reg _396909_396909 ; 
   reg __396909_396909;
   reg _396910_396910 ; 
   reg __396910_396910;
   reg _396911_396911 ; 
   reg __396911_396911;
   reg _396912_396912 ; 
   reg __396912_396912;
   reg _396913_396913 ; 
   reg __396913_396913;
   reg _396914_396914 ; 
   reg __396914_396914;
   reg _396915_396915 ; 
   reg __396915_396915;
   reg _396916_396916 ; 
   reg __396916_396916;
   reg _396917_396917 ; 
   reg __396917_396917;
   reg _396918_396918 ; 
   reg __396918_396918;
   reg _396919_396919 ; 
   reg __396919_396919;
   reg _396920_396920 ; 
   reg __396920_396920;
   reg _396921_396921 ; 
   reg __396921_396921;
   reg _396922_396922 ; 
   reg __396922_396922;
   reg _396923_396923 ; 
   reg __396923_396923;
   reg _396924_396924 ; 
   reg __396924_396924;
   reg _396925_396925 ; 
   reg __396925_396925;
   reg _396926_396926 ; 
   reg __396926_396926;
   reg _396927_396927 ; 
   reg __396927_396927;
   reg _396928_396928 ; 
   reg __396928_396928;
   reg _396929_396929 ; 
   reg __396929_396929;
   reg _396930_396930 ; 
   reg __396930_396930;
   reg _396931_396931 ; 
   reg __396931_396931;
   reg _396932_396932 ; 
   reg __396932_396932;
   reg _396933_396933 ; 
   reg __396933_396933;
   reg _396934_396934 ; 
   reg __396934_396934;
   reg _396935_396935 ; 
   reg __396935_396935;
   reg _396936_396936 ; 
   reg __396936_396936;
   reg _396937_396937 ; 
   reg __396937_396937;
   reg _396938_396938 ; 
   reg __396938_396938;
   reg _396939_396939 ; 
   reg __396939_396939;
   reg _396940_396940 ; 
   reg __396940_396940;
   reg _396941_396941 ; 
   reg __396941_396941;
   reg _396942_396942 ; 
   reg __396942_396942;
   reg _396943_396943 ; 
   reg __396943_396943;
   reg _396944_396944 ; 
   reg __396944_396944;
   reg _396945_396945 ; 
   reg __396945_396945;
   reg _396946_396946 ; 
   reg __396946_396946;
   reg _396947_396947 ; 
   reg __396947_396947;
   reg _396948_396948 ; 
   reg __396948_396948;
   reg _396949_396949 ; 
   reg __396949_396949;
   reg _396950_396950 ; 
   reg __396950_396950;
   reg _396951_396951 ; 
   reg __396951_396951;
   reg _396952_396952 ; 
   reg __396952_396952;
   reg _396953_396953 ; 
   reg __396953_396953;
   reg _396954_396954 ; 
   reg __396954_396954;
   reg _396955_396955 ; 
   reg __396955_396955;
   reg _396956_396956 ; 
   reg __396956_396956;
   reg _396957_396957 ; 
   reg __396957_396957;
   reg _396958_396958 ; 
   reg __396958_396958;
   reg _396959_396959 ; 
   reg __396959_396959;
   reg _396960_396960 ; 
   reg __396960_396960;
   reg _396961_396961 ; 
   reg __396961_396961;
   reg _396962_396962 ; 
   reg __396962_396962;
   reg _396963_396963 ; 
   reg __396963_396963;
   reg _396964_396964 ; 
   reg __396964_396964;
   reg _396965_396965 ; 
   reg __396965_396965;
   reg _396966_396966 ; 
   reg __396966_396966;
   reg _396967_396967 ; 
   reg __396967_396967;
   reg _396968_396968 ; 
   reg __396968_396968;
   reg _396969_396969 ; 
   reg __396969_396969;
   reg _396970_396970 ; 
   reg __396970_396970;
   reg _396971_396971 ; 
   reg __396971_396971;
   reg _396972_396972 ; 
   reg __396972_396972;
   reg _396973_396973 ; 
   reg __396973_396973;
   reg _396974_396974 ; 
   reg __396974_396974;
   reg _396975_396975 ; 
   reg __396975_396975;
   reg _396976_396976 ; 
   reg __396976_396976;
   reg _396977_396977 ; 
   reg __396977_396977;
   reg _396978_396978 ; 
   reg __396978_396978;
   reg _396979_396979 ; 
   reg __396979_396979;
   reg _396980_396980 ; 
   reg __396980_396980;
   reg _396981_396981 ; 
   reg __396981_396981;
   reg _396982_396982 ; 
   reg __396982_396982;
   reg _396983_396983 ; 
   reg __396983_396983;
   reg _396984_396984 ; 
   reg __396984_396984;
   reg _396985_396985 ; 
   reg __396985_396985;
   reg _396986_396986 ; 
   reg __396986_396986;
   reg _396987_396987 ; 
   reg __396987_396987;
   reg _396988_396988 ; 
   reg __396988_396988;
   reg _396989_396989 ; 
   reg __396989_396989;
   reg _396990_396990 ; 
   reg __396990_396990;
   reg _396991_396991 ; 
   reg __396991_396991;
   reg _396992_396992 ; 
   reg __396992_396992;
   reg _396993_396993 ; 
   reg __396993_396993;
   reg _396994_396994 ; 
   reg __396994_396994;
   reg _396995_396995 ; 
   reg __396995_396995;
   reg _396996_396996 ; 
   reg __396996_396996;
   reg _396997_396997 ; 
   reg __396997_396997;
   reg _396998_396998 ; 
   reg __396998_396998;
   reg _396999_396999 ; 
   reg __396999_396999;
   reg _397000_397000 ; 
   reg __397000_397000;
   reg _397001_397001 ; 
   reg __397001_397001;
   reg _397002_397002 ; 
   reg __397002_397002;
   reg _397003_397003 ; 
   reg __397003_397003;
   reg _397004_397004 ; 
   reg __397004_397004;
   reg _397005_397005 ; 
   reg __397005_397005;
   reg _397006_397006 ; 
   reg __397006_397006;
   reg _397007_397007 ; 
   reg __397007_397007;
   reg _397008_397008 ; 
   reg __397008_397008;
   reg _397009_397009 ; 
   reg __397009_397009;
   reg _397010_397010 ; 
   reg __397010_397010;
   reg _397011_397011 ; 
   reg __397011_397011;
   reg _397012_397012 ; 
   reg __397012_397012;
   reg _397013_397013 ; 
   reg __397013_397013;
   reg _397014_397014 ; 
   reg __397014_397014;
   reg _397015_397015 ; 
   reg __397015_397015;
   reg _397016_397016 ; 
   reg __397016_397016;
   reg _397017_397017 ; 
   reg __397017_397017;
   reg _397018_397018 ; 
   reg __397018_397018;
   reg _397019_397019 ; 
   reg __397019_397019;
   reg _397020_397020 ; 
   reg __397020_397020;
   reg _397021_397021 ; 
   reg __397021_397021;
   reg _397022_397022 ; 
   reg __397022_397022;
   reg _397023_397023 ; 
   reg __397023_397023;
   reg _397024_397024 ; 
   reg __397024_397024;
   reg _397025_397025 ; 
   reg __397025_397025;
   reg _397026_397026 ; 
   reg __397026_397026;
   reg _397027_397027 ; 
   reg __397027_397027;
   reg _397028_397028 ; 
   reg __397028_397028;
   reg _397029_397029 ; 
   reg __397029_397029;
   reg _397030_397030 ; 
   reg __397030_397030;
   reg _397031_397031 ; 
   reg __397031_397031;
   reg _397032_397032 ; 
   reg __397032_397032;
   reg _397033_397033 ; 
   reg __397033_397033;
   reg _397034_397034 ; 
   reg __397034_397034;
   reg _397035_397035 ; 
   reg __397035_397035;
   reg _397036_397036 ; 
   reg __397036_397036;
   reg _397037_397037 ; 
   reg __397037_397037;
   reg _397038_397038 ; 
   reg __397038_397038;
   reg _397039_397039 ; 
   reg __397039_397039;
   reg _397040_397040 ; 
   reg __397040_397040;
   reg _397041_397041 ; 
   reg __397041_397041;
   reg _397042_397042 ; 
   reg __397042_397042;
   reg _397043_397043 ; 
   reg __397043_397043;
   reg _397044_397044 ; 
   reg __397044_397044;
   reg _397045_397045 ; 
   reg __397045_397045;
   reg _397046_397046 ; 
   reg __397046_397046;
   reg _397047_397047 ; 
   reg __397047_397047;
   reg _397048_397048 ; 
   reg __397048_397048;
   reg _397049_397049 ; 
   reg __397049_397049;
   reg _397050_397050 ; 
   reg __397050_397050;
   reg _397051_397051 ; 
   reg __397051_397051;
   reg _397052_397052 ; 
   reg __397052_397052;
   reg _397053_397053 ; 
   reg __397053_397053;
   reg _397054_397054 ; 
   reg __397054_397054;
   reg _397055_397055 ; 
   reg __397055_397055;
   reg _397056_397056 ; 
   reg __397056_397056;
   reg _397057_397057 ; 
   reg __397057_397057;
   reg _397058_397058 ; 
   reg __397058_397058;
   reg _397059_397059 ; 
   reg __397059_397059;
   reg _397060_397060 ; 
   reg __397060_397060;
   reg _397061_397061 ; 
   reg __397061_397061;
   reg _397062_397062 ; 
   reg __397062_397062;
   reg _397063_397063 ; 
   reg __397063_397063;
   reg _397064_397064 ; 
   reg __397064_397064;
   reg _397065_397065 ; 
   reg __397065_397065;
   reg _397066_397066 ; 
   reg __397066_397066;
   reg _397067_397067 ; 
   reg __397067_397067;
   reg _397068_397068 ; 
   reg __397068_397068;
   reg _397069_397069 ; 
   reg __397069_397069;
   reg _397070_397070 ; 
   reg __397070_397070;
   reg _397071_397071 ; 
   reg __397071_397071;
   reg _397072_397072 ; 
   reg __397072_397072;
   reg _397073_397073 ; 
   reg __397073_397073;
   reg _397074_397074 ; 
   reg __397074_397074;
   reg _397075_397075 ; 
   reg __397075_397075;
   reg _397076_397076 ; 
   reg __397076_397076;
   reg _397077_397077 ; 
   reg __397077_397077;
   reg _397078_397078 ; 
   reg __397078_397078;
   reg _397079_397079 ; 
   reg __397079_397079;
   reg _397080_397080 ; 
   reg __397080_397080;
   reg _397081_397081 ; 
   reg __397081_397081;
   reg _397082_397082 ; 
   reg __397082_397082;
   reg _397083_397083 ; 
   reg __397083_397083;
   reg _397084_397084 ; 
   reg __397084_397084;
   reg _397085_397085 ; 
   reg __397085_397085;
   reg _397086_397086 ; 
   reg __397086_397086;
   reg _397087_397087 ; 
   reg __397087_397087;
   reg _397088_397088 ; 
   reg __397088_397088;
   reg _397089_397089 ; 
   reg __397089_397089;
   reg _397090_397090 ; 
   reg __397090_397090;
   reg _397091_397091 ; 
   reg __397091_397091;
   reg _397092_397092 ; 
   reg __397092_397092;
   reg _397093_397093 ; 
   reg __397093_397093;
   reg _397094_397094 ; 
   reg __397094_397094;
   reg _397095_397095 ; 
   reg __397095_397095;
   reg _397096_397096 ; 
   reg __397096_397096;
   reg _397097_397097 ; 
   reg __397097_397097;
   reg _397098_397098 ; 
   reg __397098_397098;
   reg _397099_397099 ; 
   reg __397099_397099;
   reg _397100_397100 ; 
   reg __397100_397100;
   reg _397101_397101 ; 
   reg __397101_397101;
   reg _397102_397102 ; 
   reg __397102_397102;
   reg _397103_397103 ; 
   reg __397103_397103;
   reg _397104_397104 ; 
   reg __397104_397104;
   reg _397105_397105 ; 
   reg __397105_397105;
   reg _397106_397106 ; 
   reg __397106_397106;
   reg _397107_397107 ; 
   reg __397107_397107;
   reg _397108_397108 ; 
   reg __397108_397108;
   reg _397109_397109 ; 
   reg __397109_397109;
   reg _397110_397110 ; 
   reg __397110_397110;
   reg _397111_397111 ; 
   reg __397111_397111;
   reg _397112_397112 ; 
   reg __397112_397112;
   reg _397113_397113 ; 
   reg __397113_397113;
   reg _397114_397114 ; 
   reg __397114_397114;
   reg _397115_397115 ; 
   reg __397115_397115;
   reg _397116_397116 ; 
   reg __397116_397116;
   reg _397117_397117 ; 
   reg __397117_397117;
   reg _397118_397118 ; 
   reg __397118_397118;
   reg _397119_397119 ; 
   reg __397119_397119;
   reg _397120_397120 ; 
   reg __397120_397120;
   reg _397121_397121 ; 
   reg __397121_397121;
   reg _397122_397122 ; 
   reg __397122_397122;
   reg _397123_397123 ; 
   reg __397123_397123;
   reg _397124_397124 ; 
   reg __397124_397124;
   reg _397125_397125 ; 
   reg __397125_397125;
   reg _397126_397126 ; 
   reg __397126_397126;
   reg _397127_397127 ; 
   reg __397127_397127;
   reg _397128_397128 ; 
   reg __397128_397128;
   reg _397129_397129 ; 
   reg __397129_397129;
   reg _397130_397130 ; 
   reg __397130_397130;
   reg _397131_397131 ; 
   reg __397131_397131;
   reg _397132_397132 ; 
   reg __397132_397132;
   reg _397133_397133 ; 
   reg __397133_397133;
   reg _397134_397134 ; 
   reg __397134_397134;
   reg _397135_397135 ; 
   reg __397135_397135;
   reg _397136_397136 ; 
   reg __397136_397136;
   reg _397137_397137 ; 
   reg __397137_397137;
   reg _397138_397138 ; 
   reg __397138_397138;
   reg _397139_397139 ; 
   reg __397139_397139;
   reg _397140_397140 ; 
   reg __397140_397140;
   reg _397141_397141 ; 
   reg __397141_397141;
   reg _397142_397142 ; 
   reg __397142_397142;
   reg _397143_397143 ; 
   reg __397143_397143;
   reg _397144_397144 ; 
   reg __397144_397144;
   reg _397145_397145 ; 
   reg __397145_397145;
   reg _397146_397146 ; 
   reg __397146_397146;
   reg _397147_397147 ; 
   reg __397147_397147;
   reg _397148_397148 ; 
   reg __397148_397148;
   reg _397149_397149 ; 
   reg __397149_397149;
   reg _397150_397150 ; 
   reg __397150_397150;
   reg _397151_397151 ; 
   reg __397151_397151;
   reg _397152_397152 ; 
   reg __397152_397152;
   reg _397153_397153 ; 
   reg __397153_397153;
   reg _397154_397154 ; 
   reg __397154_397154;
   reg _397155_397155 ; 
   reg __397155_397155;
   reg _397156_397156 ; 
   reg __397156_397156;
   reg _397157_397157 ; 
   reg __397157_397157;
   reg _397158_397158 ; 
   reg __397158_397158;
   reg _397159_397159 ; 
   reg __397159_397159;
   reg _397160_397160 ; 
   reg __397160_397160;
   reg _397161_397161 ; 
   reg __397161_397161;
   reg _397162_397162 ; 
   reg __397162_397162;
   reg _397163_397163 ; 
   reg __397163_397163;
   reg _397164_397164 ; 
   reg __397164_397164;
   reg _397165_397165 ; 
   reg __397165_397165;
   reg _397166_397166 ; 
   reg __397166_397166;
   reg _397167_397167 ; 
   reg __397167_397167;
   reg _397168_397168 ; 
   reg __397168_397168;
   reg _397169_397169 ; 
   reg __397169_397169;
   reg _397170_397170 ; 
   reg __397170_397170;
   reg _397171_397171 ; 
   reg __397171_397171;
   reg _397172_397172 ; 
   reg __397172_397172;
   reg _397173_397173 ; 
   reg __397173_397173;
   reg _397174_397174 ; 
   reg __397174_397174;
   reg _397175_397175 ; 
   reg __397175_397175;
   reg _397176_397176 ; 
   reg __397176_397176;
   reg _397177_397177 ; 
   reg __397177_397177;
   reg _397178_397178 ; 
   reg __397178_397178;
   reg _397179_397179 ; 
   reg __397179_397179;
   reg _397180_397180 ; 
   reg __397180_397180;
   reg _397181_397181 ; 
   reg __397181_397181;
   reg _397182_397182 ; 
   reg __397182_397182;
   reg _397183_397183 ; 
   reg __397183_397183;
   reg _397184_397184 ; 
   reg __397184_397184;
   reg _397185_397185 ; 
   reg __397185_397185;
   reg _397186_397186 ; 
   reg __397186_397186;
   reg _397187_397187 ; 
   reg __397187_397187;
   reg _397188_397188 ; 
   reg __397188_397188;
   reg _397189_397189 ; 
   reg __397189_397189;
   reg _397190_397190 ; 
   reg __397190_397190;
   reg _397191_397191 ; 
   reg __397191_397191;
   reg _397192_397192 ; 
   reg __397192_397192;
   reg _397193_397193 ; 
   reg __397193_397193;
   reg _397194_397194 ; 
   reg __397194_397194;
   reg _397195_397195 ; 
   reg __397195_397195;
   reg _397196_397196 ; 
   reg __397196_397196;
   reg _397197_397197 ; 
   reg __397197_397197;
   reg _397198_397198 ; 
   reg __397198_397198;
   reg _397199_397199 ; 
   reg __397199_397199;
   reg _397200_397200 ; 
   reg __397200_397200;
   reg _397201_397201 ; 
   reg __397201_397201;
   reg _397202_397202 ; 
   reg __397202_397202;
   reg _397203_397203 ; 
   reg __397203_397203;
   reg _397204_397204 ; 
   reg __397204_397204;
   reg _397205_397205 ; 
   reg __397205_397205;
   reg _397206_397206 ; 
   reg __397206_397206;
   reg _397207_397207 ; 
   reg __397207_397207;
   reg _397208_397208 ; 
   reg __397208_397208;
   reg _397209_397209 ; 
   reg __397209_397209;
   reg _397210_397210 ; 
   reg __397210_397210;
   reg _397211_397211 ; 
   reg __397211_397211;
   reg _397212_397212 ; 
   reg __397212_397212;
   reg _397213_397213 ; 
   reg __397213_397213;
   reg _397214_397214 ; 
   reg __397214_397214;
   reg _397215_397215 ; 
   reg __397215_397215;
   reg _397216_397216 ; 
   reg __397216_397216;
   reg _397217_397217 ; 
   reg __397217_397217;
   reg _397218_397218 ; 
   reg __397218_397218;
   reg _397219_397219 ; 
   reg __397219_397219;
   reg _397220_397220 ; 
   reg __397220_397220;
   reg _397221_397221 ; 
   reg __397221_397221;
   reg _397222_397222 ; 
   reg __397222_397222;
   reg _397223_397223 ; 
   reg __397223_397223;
   reg _397224_397224 ; 
   reg __397224_397224;
   reg _397225_397225 ; 
   reg __397225_397225;
   reg _397226_397226 ; 
   reg __397226_397226;
   reg _397227_397227 ; 
   reg __397227_397227;
   reg _397228_397228 ; 
   reg __397228_397228;
   reg _397229_397229 ; 
   reg __397229_397229;
   reg _397230_397230 ; 
   reg __397230_397230;
   reg _397231_397231 ; 
   reg __397231_397231;
   reg _397232_397232 ; 
   reg __397232_397232;
   reg _397233_397233 ; 
   reg __397233_397233;
   reg _397234_397234 ; 
   reg __397234_397234;
   reg _397235_397235 ; 
   reg __397235_397235;
   reg _397236_397236 ; 
   reg __397236_397236;
   reg _397237_397237 ; 
   reg __397237_397237;
   reg _397238_397238 ; 
   reg __397238_397238;
   reg _397239_397239 ; 
   reg __397239_397239;
   reg _397240_397240 ; 
   reg __397240_397240;
   reg _397241_397241 ; 
   reg __397241_397241;
   reg _397242_397242 ; 
   reg __397242_397242;
   reg _397243_397243 ; 
   reg __397243_397243;
   reg _397244_397244 ; 
   reg __397244_397244;
   reg _397245_397245 ; 
   reg __397245_397245;
   reg _397246_397246 ; 
   reg __397246_397246;
   reg _397247_397247 ; 
   reg __397247_397247;
   reg _397248_397248 ; 
   reg __397248_397248;
   reg _397249_397249 ; 
   reg __397249_397249;
   reg _397250_397250 ; 
   reg __397250_397250;
   reg _397251_397251 ; 
   reg __397251_397251;
   reg _397252_397252 ; 
   reg __397252_397252;
   reg _397253_397253 ; 
   reg __397253_397253;
   reg _397254_397254 ; 
   reg __397254_397254;
   reg _397255_397255 ; 
   reg __397255_397255;
   reg _397256_397256 ; 
   reg __397256_397256;
   reg _397257_397257 ; 
   reg __397257_397257;
   reg _397258_397258 ; 
   reg __397258_397258;
   reg _397259_397259 ; 
   reg __397259_397259;
   reg _397260_397260 ; 
   reg __397260_397260;
   reg _397261_397261 ; 
   reg __397261_397261;
   reg _397262_397262 ; 
   reg __397262_397262;
   reg _397263_397263 ; 
   reg __397263_397263;
   reg _397264_397264 ; 
   reg __397264_397264;
   reg _397265_397265 ; 
   reg __397265_397265;
   reg _397266_397266 ; 
   reg __397266_397266;
   reg _397267_397267 ; 
   reg __397267_397267;
   reg _397268_397268 ; 
   reg __397268_397268;
   reg _397269_397269 ; 
   reg __397269_397269;
   reg _397270_397270 ; 
   reg __397270_397270;
   reg _397271_397271 ; 
   reg __397271_397271;
   reg _397272_397272 ; 
   reg __397272_397272;
   reg _397273_397273 ; 
   reg __397273_397273;
   reg _397274_397274 ; 
   reg __397274_397274;
   reg _397275_397275 ; 
   reg __397275_397275;
   reg _397276_397276 ; 
   reg __397276_397276;
   reg _397277_397277 ; 
   reg __397277_397277;
   reg _397278_397278 ; 
   reg __397278_397278;
   reg _397279_397279 ; 
   reg __397279_397279;
   reg _397280_397280 ; 
   reg __397280_397280;
   reg _397281_397281 ; 
   reg __397281_397281;
   reg _397282_397282 ; 
   reg __397282_397282;
   reg _397283_397283 ; 
   reg __397283_397283;
   reg _397284_397284 ; 
   reg __397284_397284;
   reg _397285_397285 ; 
   reg __397285_397285;
   reg _397286_397286 ; 
   reg __397286_397286;
   reg _397287_397287 ; 
   reg __397287_397287;
   reg _397288_397288 ; 
   reg __397288_397288;
   reg _397289_397289 ; 
   reg __397289_397289;
   reg _397290_397290 ; 
   reg __397290_397290;
   reg _397291_397291 ; 
   reg __397291_397291;
   reg _397292_397292 ; 
   reg __397292_397292;
   reg _397293_397293 ; 
   reg __397293_397293;
   reg _397294_397294 ; 
   reg __397294_397294;
   reg _397295_397295 ; 
   reg __397295_397295;
   reg _397296_397296 ; 
   reg __397296_397296;
   reg _397297_397297 ; 
   reg __397297_397297;
   reg _397298_397298 ; 
   reg __397298_397298;
   reg _397299_397299 ; 
   reg __397299_397299;
   reg _397300_397300 ; 
   reg __397300_397300;
   reg _397301_397301 ; 
   reg __397301_397301;
   reg _397302_397302 ; 
   reg __397302_397302;
   reg _397303_397303 ; 
   reg __397303_397303;
   reg _397304_397304 ; 
   reg __397304_397304;
   reg _397305_397305 ; 
   reg __397305_397305;
   reg _397306_397306 ; 
   reg __397306_397306;
   reg _397307_397307 ; 
   reg __397307_397307;
   reg _397308_397308 ; 
   reg __397308_397308;
   reg _397309_397309 ; 
   reg __397309_397309;
   reg _397310_397310 ; 
   reg __397310_397310;
   reg _397311_397311 ; 
   reg __397311_397311;
   reg _397312_397312 ; 
   reg __397312_397312;
   reg _397313_397313 ; 
   reg __397313_397313;
   reg _397314_397314 ; 
   reg __397314_397314;
   reg _397315_397315 ; 
   reg __397315_397315;
   reg _397316_397316 ; 
   reg __397316_397316;
   reg _397317_397317 ; 
   reg __397317_397317;
   reg _397318_397318 ; 
   reg __397318_397318;
   reg _397319_397319 ; 
   reg __397319_397319;
   reg _397320_397320 ; 
   reg __397320_397320;
   reg _397321_397321 ; 
   reg __397321_397321;
   reg _397322_397322 ; 
   reg __397322_397322;
   reg _397323_397323 ; 
   reg __397323_397323;
   reg _397324_397324 ; 
   reg __397324_397324;
   reg _397325_397325 ; 
   reg __397325_397325;
   reg _397326_397326 ; 
   reg __397326_397326;
   reg _397327_397327 ; 
   reg __397327_397327;
   reg _397328_397328 ; 
   reg __397328_397328;
   reg _397329_397329 ; 
   reg __397329_397329;
   reg _397330_397330 ; 
   reg __397330_397330;
   reg _397331_397331 ; 
   reg __397331_397331;
   reg _397332_397332 ; 
   reg __397332_397332;
   reg _397333_397333 ; 
   reg __397333_397333;
   reg _397334_397334 ; 
   reg __397334_397334;
   reg _397335_397335 ; 
   reg __397335_397335;
   reg _397336_397336 ; 
   reg __397336_397336;
   reg _397337_397337 ; 
   reg __397337_397337;
   reg _397338_397338 ; 
   reg __397338_397338;
   reg _397339_397339 ; 
   reg __397339_397339;
   reg _397340_397340 ; 
   reg __397340_397340;
   reg _397341_397341 ; 
   reg __397341_397341;
   reg _397342_397342 ; 
   reg __397342_397342;
   reg _397343_397343 ; 
   reg __397343_397343;
   reg _397344_397344 ; 
   reg __397344_397344;
   reg _397345_397345 ; 
   reg __397345_397345;
   reg _397346_397346 ; 
   reg __397346_397346;
   reg _397347_397347 ; 
   reg __397347_397347;
   reg _397348_397348 ; 
   reg __397348_397348;
   reg _397349_397349 ; 
   reg __397349_397349;
   reg _397350_397350 ; 
   reg __397350_397350;
   reg _397351_397351 ; 
   reg __397351_397351;
   reg _397352_397352 ; 
   reg __397352_397352;
   reg _397353_397353 ; 
   reg __397353_397353;
   reg _397354_397354 ; 
   reg __397354_397354;
   reg _397355_397355 ; 
   reg __397355_397355;
   reg _397356_397356 ; 
   reg __397356_397356;
   reg _397357_397357 ; 
   reg __397357_397357;
   reg _397358_397358 ; 
   reg __397358_397358;
   reg _397359_397359 ; 
   reg __397359_397359;
   reg _397360_397360 ; 
   reg __397360_397360;
   reg _397361_397361 ; 
   reg __397361_397361;
   reg _397362_397362 ; 
   reg __397362_397362;
   reg _397363_397363 ; 
   reg __397363_397363;
   reg _397364_397364 ; 
   reg __397364_397364;
   reg _397365_397365 ; 
   reg __397365_397365;
   reg _397366_397366 ; 
   reg __397366_397366;
   reg _397367_397367 ; 
   reg __397367_397367;
   reg _397368_397368 ; 
   reg __397368_397368;
   reg _397369_397369 ; 
   reg __397369_397369;
   reg _397370_397370 ; 
   reg __397370_397370;
   reg _397371_397371 ; 
   reg __397371_397371;
   reg _397372_397372 ; 
   reg __397372_397372;
   reg _397373_397373 ; 
   reg __397373_397373;
   reg _397374_397374 ; 
   reg __397374_397374;
   reg _397375_397375 ; 
   reg __397375_397375;
   reg _397376_397376 ; 
   reg __397376_397376;
   reg _397377_397377 ; 
   reg __397377_397377;
   reg _397378_397378 ; 
   reg __397378_397378;
   reg _397379_397379 ; 
   reg __397379_397379;
   reg _397380_397380 ; 
   reg __397380_397380;
   reg _397381_397381 ; 
   reg __397381_397381;
   reg _397382_397382 ; 
   reg __397382_397382;
   reg _397383_397383 ; 
   reg __397383_397383;
   reg _397384_397384 ; 
   reg __397384_397384;
   reg _397385_397385 ; 
   reg __397385_397385;
   reg _397386_397386 ; 
   reg __397386_397386;
   reg _397387_397387 ; 
   reg __397387_397387;
   reg _397388_397388 ; 
   reg __397388_397388;
   reg _397389_397389 ; 
   reg __397389_397389;
   reg _397390_397390 ; 
   reg __397390_397390;
   reg _397391_397391 ; 
   reg __397391_397391;
   reg _397392_397392 ; 
   reg __397392_397392;
   reg _397393_397393 ; 
   reg __397393_397393;
   reg _397394_397394 ; 
   reg __397394_397394;
   reg _397395_397395 ; 
   reg __397395_397395;
   reg _397396_397396 ; 
   reg __397396_397396;
   reg _397397_397397 ; 
   reg __397397_397397;
   reg _397398_397398 ; 
   reg __397398_397398;
   reg _397399_397399 ; 
   reg __397399_397399;
   reg _397400_397400 ; 
   reg __397400_397400;
   reg _397401_397401 ; 
   reg __397401_397401;
   reg _397402_397402 ; 
   reg __397402_397402;
   reg _397403_397403 ; 
   reg __397403_397403;
   reg _397404_397404 ; 
   reg __397404_397404;
   reg _397405_397405 ; 
   reg __397405_397405;
   reg _397406_397406 ; 
   reg __397406_397406;
   reg _397407_397407 ; 
   reg __397407_397407;
   reg _397408_397408 ; 
   reg __397408_397408;
   reg _397409_397409 ; 
   reg __397409_397409;
   reg _397410_397410 ; 
   reg __397410_397410;
   reg _397411_397411 ; 
   reg __397411_397411;
   reg _397412_397412 ; 
   reg __397412_397412;
   reg _397413_397413 ; 
   reg __397413_397413;
   reg _397414_397414 ; 
   reg __397414_397414;
   reg _397415_397415 ; 
   reg __397415_397415;
   reg _397416_397416 ; 
   reg __397416_397416;
   reg _397417_397417 ; 
   reg __397417_397417;
   reg _397418_397418 ; 
   reg __397418_397418;
   reg _397419_397419 ; 
   reg __397419_397419;
   reg _397420_397420 ; 
   reg __397420_397420;
   reg _397421_397421 ; 
   reg __397421_397421;
   reg _397422_397422 ; 
   reg __397422_397422;
   reg _397423_397423 ; 
   reg __397423_397423;
   reg _397424_397424 ; 
   reg __397424_397424;
   reg _397425_397425 ; 
   reg __397425_397425;
   reg _397426_397426 ; 
   reg __397426_397426;
   reg _397427_397427 ; 
   reg __397427_397427;
   reg _397428_397428 ; 
   reg __397428_397428;
   reg _397429_397429 ; 
   reg __397429_397429;
   reg _397430_397430 ; 
   reg __397430_397430;
   reg _397431_397431 ; 
   reg __397431_397431;
   reg _397432_397432 ; 
   reg __397432_397432;
   reg _397433_397433 ; 
   reg __397433_397433;
   reg _397434_397434 ; 
   reg __397434_397434;
   reg _397435_397435 ; 
   reg __397435_397435;
   reg _397436_397436 ; 
   reg __397436_397436;
   reg _397437_397437 ; 
   reg __397437_397437;
   reg _397438_397438 ; 
   reg __397438_397438;
   reg _397439_397439 ; 
   reg __397439_397439;
   reg _397440_397440 ; 
   reg __397440_397440;
   reg _397441_397441 ; 
   reg __397441_397441;
   reg _397442_397442 ; 
   reg __397442_397442;
   reg _397443_397443 ; 
   reg __397443_397443;
   reg _397444_397444 ; 
   reg __397444_397444;
   reg _397445_397445 ; 
   reg __397445_397445;
   reg _397446_397446 ; 
   reg __397446_397446;
   reg _397447_397447 ; 
   reg __397447_397447;
   reg _397448_397448 ; 
   reg __397448_397448;
   reg _397449_397449 ; 
   reg __397449_397449;
   reg _397450_397450 ; 
   reg __397450_397450;
   reg _397451_397451 ; 
   reg __397451_397451;
   reg _397452_397452 ; 
   reg __397452_397452;
   reg _397453_397453 ; 
   reg __397453_397453;
   reg _397454_397454 ; 
   reg __397454_397454;
   reg _397455_397455 ; 
   reg __397455_397455;
   reg _397456_397456 ; 
   reg __397456_397456;
   reg _397457_397457 ; 
   reg __397457_397457;
   reg _397458_397458 ; 
   reg __397458_397458;
   reg _397459_397459 ; 
   reg __397459_397459;
   reg _397460_397460 ; 
   reg __397460_397460;
   reg _397461_397461 ; 
   reg __397461_397461;
   reg _397462_397462 ; 
   reg __397462_397462;
   reg _397463_397463 ; 
   reg __397463_397463;
   reg _397464_397464 ; 
   reg __397464_397464;
   reg _397465_397465 ; 
   reg __397465_397465;
   reg _397466_397466 ; 
   reg __397466_397466;
   reg _397467_397467 ; 
   reg __397467_397467;
   reg _397468_397468 ; 
   reg __397468_397468;
   reg _397469_397469 ; 
   reg __397469_397469;
   reg _397470_397470 ; 
   reg __397470_397470;
   reg _397471_397471 ; 
   reg __397471_397471;
   reg _397472_397472 ; 
   reg __397472_397472;
   reg _397473_397473 ; 
   reg __397473_397473;
   reg _397474_397474 ; 
   reg __397474_397474;
   reg _397475_397475 ; 
   reg __397475_397475;
   reg _397476_397476 ; 
   reg __397476_397476;
   reg _397477_397477 ; 
   reg __397477_397477;
   reg _397478_397478 ; 
   reg __397478_397478;
   reg _397479_397479 ; 
   reg __397479_397479;
   reg _397480_397480 ; 
   reg __397480_397480;
   reg _397481_397481 ; 
   reg __397481_397481;
   reg _397482_397482 ; 
   reg __397482_397482;
   reg _397483_397483 ; 
   reg __397483_397483;
   reg _397484_397484 ; 
   reg __397484_397484;
   reg _397485_397485 ; 
   reg __397485_397485;
   reg _397486_397486 ; 
   reg __397486_397486;
   reg _397487_397487 ; 
   reg __397487_397487;
   reg _397488_397488 ; 
   reg __397488_397488;
   reg _397489_397489 ; 
   reg __397489_397489;
   reg _397490_397490 ; 
   reg __397490_397490;
   reg _397491_397491 ; 
   reg __397491_397491;
   reg _397492_397492 ; 
   reg __397492_397492;
   reg _397493_397493 ; 
   reg __397493_397493;
   reg _397494_397494 ; 
   reg __397494_397494;
   reg _397495_397495 ; 
   reg __397495_397495;
   reg _397496_397496 ; 
   reg __397496_397496;
   reg _397497_397497 ; 
   reg __397497_397497;
   reg _397498_397498 ; 
   reg __397498_397498;
   reg _397499_397499 ; 
   reg __397499_397499;
   reg _397500_397500 ; 
   reg __397500_397500;
   reg _397501_397501 ; 
   reg __397501_397501;
   reg _397502_397502 ; 
   reg __397502_397502;
   reg _397503_397503 ; 
   reg __397503_397503;
   reg _397504_397504 ; 
   reg __397504_397504;
   reg _397505_397505 ; 
   reg __397505_397505;
   reg _397506_397506 ; 
   reg __397506_397506;
   reg _397507_397507 ; 
   reg __397507_397507;
   reg _397508_397508 ; 
   reg __397508_397508;
   reg _397509_397509 ; 
   reg __397509_397509;
   reg _397510_397510 ; 
   reg __397510_397510;
   reg _397511_397511 ; 
   reg __397511_397511;
   reg _397512_397512 ; 
   reg __397512_397512;
   reg _397513_397513 ; 
   reg __397513_397513;
   reg _397514_397514 ; 
   reg __397514_397514;
   reg _397515_397515 ; 
   reg __397515_397515;
   reg _397516_397516 ; 
   reg __397516_397516;
   reg _397517_397517 ; 
   reg __397517_397517;
   reg _397518_397518 ; 
   reg __397518_397518;
   reg _397519_397519 ; 
   reg __397519_397519;
   reg _397520_397520 ; 
   reg __397520_397520;
   reg _397521_397521 ; 
   reg __397521_397521;
   reg _397522_397522 ; 
   reg __397522_397522;
   reg _397523_397523 ; 
   reg __397523_397523;
   reg _397524_397524 ; 
   reg __397524_397524;
   reg _397525_397525 ; 
   reg __397525_397525;
   reg _397526_397526 ; 
   reg __397526_397526;
   reg _397527_397527 ; 
   reg __397527_397527;
   reg _397528_397528 ; 
   reg __397528_397528;
   reg _397529_397529 ; 
   reg __397529_397529;
   reg _397530_397530 ; 
   reg __397530_397530;
   reg _397531_397531 ; 
   reg __397531_397531;
   reg _397532_397532 ; 
   reg __397532_397532;
   reg _397533_397533 ; 
   reg __397533_397533;
   reg _397534_397534 ; 
   reg __397534_397534;
   reg _397535_397535 ; 
   reg __397535_397535;
   reg _397536_397536 ; 
   reg __397536_397536;
   reg _397537_397537 ; 
   reg __397537_397537;
   reg _397538_397538 ; 
   reg __397538_397538;
   reg _397539_397539 ; 
   reg __397539_397539;
   reg _397540_397540 ; 
   reg __397540_397540;
   reg _397541_397541 ; 
   reg __397541_397541;
   reg _397542_397542 ; 
   reg __397542_397542;
   reg _397543_397543 ; 
   reg __397543_397543;
   reg _397544_397544 ; 
   reg __397544_397544;
   reg _397545_397545 ; 
   reg __397545_397545;
   reg _397546_397546 ; 
   reg __397546_397546;
   reg _397547_397547 ; 
   reg __397547_397547;
   reg _397548_397548 ; 
   reg __397548_397548;
   reg _397549_397549 ; 
   reg __397549_397549;
   reg _397550_397550 ; 
   reg __397550_397550;
   reg _397551_397551 ; 
   reg __397551_397551;
   reg _397552_397552 ; 
   reg __397552_397552;
   reg _397553_397553 ; 
   reg __397553_397553;
   reg _397554_397554 ; 
   reg __397554_397554;
   reg _397555_397555 ; 
   reg __397555_397555;
   reg _397556_397556 ; 
   reg __397556_397556;
   reg _397557_397557 ; 
   reg __397557_397557;
   reg _397558_397558 ; 
   reg __397558_397558;
   reg _397559_397559 ; 
   reg __397559_397559;
   reg _397560_397560 ; 
   reg __397560_397560;
   reg _397561_397561 ; 
   reg __397561_397561;
   reg _397562_397562 ; 
   reg __397562_397562;
   reg _397563_397563 ; 
   reg __397563_397563;
   reg _397564_397564 ; 
   reg __397564_397564;
   reg _397565_397565 ; 
   reg __397565_397565;
   reg _397566_397566 ; 
   reg __397566_397566;
   reg _397567_397567 ; 
   reg __397567_397567;
   reg _397568_397568 ; 
   reg __397568_397568;
   reg _397569_397569 ; 
   reg __397569_397569;
   reg _397570_397570 ; 
   reg __397570_397570;
   reg _397571_397571 ; 
   reg __397571_397571;
   reg _397572_397572 ; 
   reg __397572_397572;
   reg _397573_397573 ; 
   reg __397573_397573;
   reg _397574_397574 ; 
   reg __397574_397574;
   reg _397575_397575 ; 
   reg __397575_397575;
   reg _397576_397576 ; 
   reg __397576_397576;
   reg _397577_397577 ; 
   reg __397577_397577;
   reg _397578_397578 ; 
   reg __397578_397578;
   reg _397579_397579 ; 
   reg __397579_397579;
   reg _397580_397580 ; 
   reg __397580_397580;
   reg _397581_397581 ; 
   reg __397581_397581;
   reg _397582_397582 ; 
   reg __397582_397582;
   reg _397583_397583 ; 
   reg __397583_397583;
   reg _397584_397584 ; 
   reg __397584_397584;
   reg _397585_397585 ; 
   reg __397585_397585;
   reg _397586_397586 ; 
   reg __397586_397586;
   reg _397587_397587 ; 
   reg __397587_397587;
   reg _397588_397588 ; 
   reg __397588_397588;
   reg _397589_397589 ; 
   reg __397589_397589;
   reg _397590_397590 ; 
   reg __397590_397590;
   reg _397591_397591 ; 
   reg __397591_397591;
   reg _397592_397592 ; 
   reg __397592_397592;
   reg _397593_397593 ; 
   reg __397593_397593;
   reg _397594_397594 ; 
   reg __397594_397594;
   reg _397595_397595 ; 
   reg __397595_397595;
   reg _397596_397596 ; 
   reg __397596_397596;
   reg _397597_397597 ; 
   reg __397597_397597;
   reg _397598_397598 ; 
   reg __397598_397598;
   reg _397599_397599 ; 
   reg __397599_397599;
   reg _397600_397600 ; 
   reg __397600_397600;
   reg _397601_397601 ; 
   reg __397601_397601;
   reg _397602_397602 ; 
   reg __397602_397602;
   reg _397603_397603 ; 
   reg __397603_397603;
   reg _397604_397604 ; 
   reg __397604_397604;
   reg _397605_397605 ; 
   reg __397605_397605;
   reg _397606_397606 ; 
   reg __397606_397606;
   reg _397607_397607 ; 
   reg __397607_397607;
   reg _397608_397608 ; 
   reg __397608_397608;
   reg _397609_397609 ; 
   reg __397609_397609;
   reg _397610_397610 ; 
   reg __397610_397610;
   reg _397611_397611 ; 
   reg __397611_397611;
   reg _397612_397612 ; 
   reg __397612_397612;
   reg _397613_397613 ; 
   reg __397613_397613;
   reg _397614_397614 ; 
   reg __397614_397614;
   reg _397615_397615 ; 
   reg __397615_397615;
   reg _397616_397616 ; 
   reg __397616_397616;
   reg _397617_397617 ; 
   reg __397617_397617;
   reg _397618_397618 ; 
   reg __397618_397618;
   reg _397619_397619 ; 
   reg __397619_397619;
   reg _397620_397620 ; 
   reg __397620_397620;
   reg _397621_397621 ; 
   reg __397621_397621;
   reg _397622_397622 ; 
   reg __397622_397622;
   reg _397623_397623 ; 
   reg __397623_397623;
   reg _397624_397624 ; 
   reg __397624_397624;
   reg _397625_397625 ; 
   reg __397625_397625;
   reg _397626_397626 ; 
   reg __397626_397626;
   reg _397627_397627 ; 
   reg __397627_397627;
   reg _397628_397628 ; 
   reg __397628_397628;
   reg _397629_397629 ; 
   reg __397629_397629;
   reg _397630_397630 ; 
   reg __397630_397630;
   reg _397631_397631 ; 
   reg __397631_397631;
   reg _397632_397632 ; 
   reg __397632_397632;
   reg _397633_397633 ; 
   reg __397633_397633;
   reg _397634_397634 ; 
   reg __397634_397634;
   reg _397635_397635 ; 
   reg __397635_397635;
   reg _397636_397636 ; 
   reg __397636_397636;
   reg _397637_397637 ; 
   reg __397637_397637;
   reg _397638_397638 ; 
   reg __397638_397638;
   reg _397639_397639 ; 
   reg __397639_397639;
   reg _397640_397640 ; 
   reg __397640_397640;
   reg _397641_397641 ; 
   reg __397641_397641;
   reg _397642_397642 ; 
   reg __397642_397642;
   reg _397643_397643 ; 
   reg __397643_397643;
   reg _397644_397644 ; 
   reg __397644_397644;
   reg _397645_397645 ; 
   reg __397645_397645;
   reg _397646_397646 ; 
   reg __397646_397646;
   reg _397647_397647 ; 
   reg __397647_397647;
   reg _397648_397648 ; 
   reg __397648_397648;
   reg _397649_397649 ; 
   reg __397649_397649;
   reg _397650_397650 ; 
   reg __397650_397650;
   reg _397651_397651 ; 
   reg __397651_397651;
   reg _397652_397652 ; 
   reg __397652_397652;
   reg _397653_397653 ; 
   reg __397653_397653;
   reg _397654_397654 ; 
   reg __397654_397654;
   reg _397655_397655 ; 
   reg __397655_397655;
   reg _397656_397656 ; 
   reg __397656_397656;
   reg _397657_397657 ; 
   reg __397657_397657;
   reg _397658_397658 ; 
   reg __397658_397658;
   reg _397659_397659 ; 
   reg __397659_397659;
   reg _397660_397660 ; 
   reg __397660_397660;
   reg _397661_397661 ; 
   reg __397661_397661;
   reg _397662_397662 ; 
   reg __397662_397662;
   reg _397663_397663 ; 
   reg __397663_397663;
   reg _397664_397664 ; 
   reg __397664_397664;
   reg _397665_397665 ; 
   reg __397665_397665;
   reg _397666_397666 ; 
   reg __397666_397666;
   reg _397667_397667 ; 
   reg __397667_397667;
   reg _397668_397668 ; 
   reg __397668_397668;
   reg _397669_397669 ; 
   reg __397669_397669;
   reg _397670_397670 ; 
   reg __397670_397670;
   reg _397671_397671 ; 
   reg __397671_397671;
   reg _397672_397672 ; 
   reg __397672_397672;
   reg _397673_397673 ; 
   reg __397673_397673;
   reg _397674_397674 ; 
   reg __397674_397674;
   reg _397675_397675 ; 
   reg __397675_397675;
   reg _397676_397676 ; 
   reg __397676_397676;
   reg _397677_397677 ; 
   reg __397677_397677;
   reg _397678_397678 ; 
   reg __397678_397678;
   reg _397679_397679 ; 
   reg __397679_397679;
   reg _397680_397680 ; 
   reg __397680_397680;
   reg _397681_397681 ; 
   reg __397681_397681;
   reg _397682_397682 ; 
   reg __397682_397682;
   reg _397683_397683 ; 
   reg __397683_397683;
   reg _397684_397684 ; 
   reg __397684_397684;
   reg _397685_397685 ; 
   reg __397685_397685;
   reg _397686_397686 ; 
   reg __397686_397686;
   reg _397687_397687 ; 
   reg __397687_397687;
   reg _397688_397688 ; 
   reg __397688_397688;
   reg _397689_397689 ; 
   reg __397689_397689;
   reg _397690_397690 ; 
   reg __397690_397690;
   reg _397691_397691 ; 
   reg __397691_397691;
   reg _397692_397692 ; 
   reg __397692_397692;
   reg _397693_397693 ; 
   reg __397693_397693;
   reg _397694_397694 ; 
   reg __397694_397694;
   reg _397695_397695 ; 
   reg __397695_397695;
   reg _397696_397696 ; 
   reg __397696_397696;
   reg _397697_397697 ; 
   reg __397697_397697;
   reg _397698_397698 ; 
   reg __397698_397698;
   reg _397699_397699 ; 
   reg __397699_397699;
   reg _397700_397700 ; 
   reg __397700_397700;
   reg _397701_397701 ; 
   reg __397701_397701;
   reg _397702_397702 ; 
   reg __397702_397702;
   reg _397703_397703 ; 
   reg __397703_397703;
   reg _397704_397704 ; 
   reg __397704_397704;
   reg _397705_397705 ; 
   reg __397705_397705;
   reg _397706_397706 ; 
   reg __397706_397706;
   reg _397707_397707 ; 
   reg __397707_397707;
   reg _397708_397708 ; 
   reg __397708_397708;
   reg _397709_397709 ; 
   reg __397709_397709;
   reg _397710_397710 ; 
   reg __397710_397710;
   reg _397711_397711 ; 
   reg __397711_397711;
   reg _397712_397712 ; 
   reg __397712_397712;
   reg _397713_397713 ; 
   reg __397713_397713;
   reg _397714_397714 ; 
   reg __397714_397714;
   reg _397715_397715 ; 
   reg __397715_397715;
   reg _397716_397716 ; 
   reg __397716_397716;
   reg _397717_397717 ; 
   reg __397717_397717;
   reg _397718_397718 ; 
   reg __397718_397718;
   reg _397719_397719 ; 
   reg __397719_397719;
   reg _397720_397720 ; 
   reg __397720_397720;
   reg _397721_397721 ; 
   reg __397721_397721;
   reg _397722_397722 ; 
   reg __397722_397722;
   reg _397723_397723 ; 
   reg __397723_397723;
   reg _397724_397724 ; 
   reg __397724_397724;
   reg _397725_397725 ; 
   reg __397725_397725;
   reg _397726_397726 ; 
   reg __397726_397726;
   reg _397727_397727 ; 
   reg __397727_397727;
   reg _397728_397728 ; 
   reg __397728_397728;
   reg _397729_397729 ; 
   reg __397729_397729;
   reg _397730_397730 ; 
   reg __397730_397730;
   reg _397731_397731 ; 
   reg __397731_397731;
   reg _397732_397732 ; 
   reg __397732_397732;
   reg _397733_397733 ; 
   reg __397733_397733;
   reg _397734_397734 ; 
   reg __397734_397734;
   reg _397735_397735 ; 
   reg __397735_397735;
   reg _397736_397736 ; 
   reg __397736_397736;
   reg _397737_397737 ; 
   reg __397737_397737;
   reg _397738_397738 ; 
   reg __397738_397738;
   reg _397739_397739 ; 
   reg __397739_397739;
   reg _397740_397740 ; 
   reg __397740_397740;
   reg _397741_397741 ; 
   reg __397741_397741;
   reg _397742_397742 ; 
   reg __397742_397742;
   reg _397743_397743 ; 
   reg __397743_397743;
   reg _397744_397744 ; 
   reg __397744_397744;
   reg _397745_397745 ; 
   reg __397745_397745;
   reg _397746_397746 ; 
   reg __397746_397746;
   reg _397747_397747 ; 
   reg __397747_397747;
   reg _397748_397748 ; 
   reg __397748_397748;
   reg _397749_397749 ; 
   reg __397749_397749;
   reg _397750_397750 ; 
   reg __397750_397750;
   reg _397751_397751 ; 
   reg __397751_397751;
   reg _397752_397752 ; 
   reg __397752_397752;
   reg _397753_397753 ; 
   reg __397753_397753;
   reg _397754_397754 ; 
   reg __397754_397754;
   reg _397755_397755 ; 
   reg __397755_397755;
   reg _397756_397756 ; 
   reg __397756_397756;
   reg _397757_397757 ; 
   reg __397757_397757;
   reg _397758_397758 ; 
   reg __397758_397758;
   reg _397759_397759 ; 
   reg __397759_397759;
   reg _397760_397760 ; 
   reg __397760_397760;
   reg _397761_397761 ; 
   reg __397761_397761;
   reg _397762_397762 ; 
   reg __397762_397762;
   reg _397763_397763 ; 
   reg __397763_397763;
   reg _397764_397764 ; 
   reg __397764_397764;
   reg _397765_397765 ; 
   reg __397765_397765;
   reg _397766_397766 ; 
   reg __397766_397766;
   reg _397767_397767 ; 
   reg __397767_397767;
   reg _397768_397768 ; 
   reg __397768_397768;
   reg _397769_397769 ; 
   reg __397769_397769;
   reg _397770_397770 ; 
   reg __397770_397770;
   reg _397771_397771 ; 
   reg __397771_397771;
   reg _397772_397772 ; 
   reg __397772_397772;
   reg _397773_397773 ; 
   reg __397773_397773;
   reg _397774_397774 ; 
   reg __397774_397774;
   reg _397775_397775 ; 
   reg __397775_397775;
   reg _397776_397776 ; 
   reg __397776_397776;
   reg _397777_397777 ; 
   reg __397777_397777;
   reg _397778_397778 ; 
   reg __397778_397778;
   reg _397779_397779 ; 
   reg __397779_397779;
   reg _397780_397780 ; 
   reg __397780_397780;
   reg _397781_397781 ; 
   reg __397781_397781;
   reg _397782_397782 ; 
   reg __397782_397782;
   reg _397783_397783 ; 
   reg __397783_397783;
   reg _397784_397784 ; 
   reg __397784_397784;
   reg _397785_397785 ; 
   reg __397785_397785;
   reg _397786_397786 ; 
   reg __397786_397786;
   reg _397787_397787 ; 
   reg __397787_397787;
   reg _397788_397788 ; 
   reg __397788_397788;
   reg _397789_397789 ; 
   reg __397789_397789;
   reg _397790_397790 ; 
   reg __397790_397790;
   reg _397791_397791 ; 
   reg __397791_397791;
   reg _397792_397792 ; 
   reg __397792_397792;
   reg _397793_397793 ; 
   reg __397793_397793;
   reg _397794_397794 ; 
   reg __397794_397794;
   reg _397795_397795 ; 
   reg __397795_397795;
   reg _397796_397796 ; 
   reg __397796_397796;
   reg _397797_397797 ; 
   reg __397797_397797;
   reg _397798_397798 ; 
   reg __397798_397798;
   reg _397799_397799 ; 
   reg __397799_397799;
   reg _397800_397800 ; 
   reg __397800_397800;
   reg _397801_397801 ; 
   reg __397801_397801;
   reg _397802_397802 ; 
   reg __397802_397802;
   reg _397803_397803 ; 
   reg __397803_397803;
   reg _397804_397804 ; 
   reg __397804_397804;
   reg _397805_397805 ; 
   reg __397805_397805;
   reg _397806_397806 ; 
   reg __397806_397806;
   reg _397807_397807 ; 
   reg __397807_397807;
   reg _397808_397808 ; 
   reg __397808_397808;
   reg _397809_397809 ; 
   reg __397809_397809;
   reg _397810_397810 ; 
   reg __397810_397810;
   reg _397811_397811 ; 
   reg __397811_397811;
   reg _397812_397812 ; 
   reg __397812_397812;
   reg _397813_397813 ; 
   reg __397813_397813;
   reg _397814_397814 ; 
   reg __397814_397814;
   reg _397815_397815 ; 
   reg __397815_397815;
   reg _397816_397816 ; 
   reg __397816_397816;
   reg _397817_397817 ; 
   reg __397817_397817;
   reg _397818_397818 ; 
   reg __397818_397818;
   reg _397819_397819 ; 
   reg __397819_397819;
   reg _397820_397820 ; 
   reg __397820_397820;
   reg _397821_397821 ; 
   reg __397821_397821;
   reg _397822_397822 ; 
   reg __397822_397822;
   reg _397823_397823 ; 
   reg __397823_397823;
   reg _397824_397824 ; 
   reg __397824_397824;
   reg _397825_397825 ; 
   reg __397825_397825;
   reg _397826_397826 ; 
   reg __397826_397826;
   reg _397827_397827 ; 
   reg __397827_397827;
   reg _397828_397828 ; 
   reg __397828_397828;
   reg _397829_397829 ; 
   reg __397829_397829;
   reg _397830_397830 ; 
   reg __397830_397830;
   reg _397831_397831 ; 
   reg __397831_397831;
   reg _397832_397832 ; 
   reg __397832_397832;
   reg _397833_397833 ; 
   reg __397833_397833;
   reg _397834_397834 ; 
   reg __397834_397834;
   reg _397835_397835 ; 
   reg __397835_397835;
   reg _397836_397836 ; 
   reg __397836_397836;
   reg _397837_397837 ; 
   reg __397837_397837;
   reg _397838_397838 ; 
   reg __397838_397838;
   reg _397839_397839 ; 
   reg __397839_397839;
   reg _397840_397840 ; 
   reg __397840_397840;
   reg _397841_397841 ; 
   reg __397841_397841;
   reg _397842_397842 ; 
   reg __397842_397842;
   reg _397843_397843 ; 
   reg __397843_397843;
   reg _397844_397844 ; 
   reg __397844_397844;
   reg _397845_397845 ; 
   reg __397845_397845;
   reg _397846_397846 ; 
   reg __397846_397846;
   reg _397847_397847 ; 
   reg __397847_397847;
   reg _397848_397848 ; 
   reg __397848_397848;
   reg _397849_397849 ; 
   reg __397849_397849;
   reg _397850_397850 ; 
   reg __397850_397850;
   reg _397851_397851 ; 
   reg __397851_397851;
   reg _397852_397852 ; 
   reg __397852_397852;
   reg _397853_397853 ; 
   reg __397853_397853;
   reg _397854_397854 ; 
   reg __397854_397854;
   reg _397855_397855 ; 
   reg __397855_397855;
   reg _397856_397856 ; 
   reg __397856_397856;
   reg _397857_397857 ; 
   reg __397857_397857;
   reg _397858_397858 ; 
   reg __397858_397858;
   reg _397859_397859 ; 
   reg __397859_397859;
   reg _397860_397860 ; 
   reg __397860_397860;
   reg _397861_397861 ; 
   reg __397861_397861;
   reg _397862_397862 ; 
   reg __397862_397862;
   reg _397863_397863 ; 
   reg __397863_397863;
   reg _397864_397864 ; 
   reg __397864_397864;
   reg _397865_397865 ; 
   reg __397865_397865;
   reg _397866_397866 ; 
   reg __397866_397866;
   reg _397867_397867 ; 
   reg __397867_397867;
   reg _397868_397868 ; 
   reg __397868_397868;
   reg _397869_397869 ; 
   reg __397869_397869;
   reg _397870_397870 ; 
   reg __397870_397870;
   reg _397871_397871 ; 
   reg __397871_397871;
   reg _397872_397872 ; 
   reg __397872_397872;
   reg _397873_397873 ; 
   reg __397873_397873;
   reg _397874_397874 ; 
   reg __397874_397874;
   reg _397875_397875 ; 
   reg __397875_397875;
   reg _397876_397876 ; 
   reg __397876_397876;
   reg _397877_397877 ; 
   reg __397877_397877;
   reg _397878_397878 ; 
   reg __397878_397878;
   reg _397879_397879 ; 
   reg __397879_397879;
   reg _397880_397880 ; 
   reg __397880_397880;
   reg _397881_397881 ; 
   reg __397881_397881;
   reg _397882_397882 ; 
   reg __397882_397882;
   reg _397883_397883 ; 
   reg __397883_397883;
   reg _397884_397884 ; 
   reg __397884_397884;
   reg _397885_397885 ; 
   reg __397885_397885;
   reg _397886_397886 ; 
   reg __397886_397886;
   reg _397887_397887 ; 
   reg __397887_397887;
   reg _397888_397888 ; 
   reg __397888_397888;
   reg _397889_397889 ; 
   reg __397889_397889;
   reg _397890_397890 ; 
   reg __397890_397890;
   reg _397891_397891 ; 
   reg __397891_397891;
   reg _397892_397892 ; 
   reg __397892_397892;
   reg _397893_397893 ; 
   reg __397893_397893;
   reg _397894_397894 ; 
   reg __397894_397894;
   reg _397895_397895 ; 
   reg __397895_397895;
   reg _397896_397896 ; 
   reg __397896_397896;
   reg _397897_397897 ; 
   reg __397897_397897;
   reg _397898_397898 ; 
   reg __397898_397898;
   reg _397899_397899 ; 
   reg __397899_397899;
   reg _397900_397900 ; 
   reg __397900_397900;
   reg _397901_397901 ; 
   reg __397901_397901;
   reg _397902_397902 ; 
   reg __397902_397902;
   reg _397903_397903 ; 
   reg __397903_397903;
   reg _397904_397904 ; 
   reg __397904_397904;
   reg _397905_397905 ; 
   reg __397905_397905;
   reg _397906_397906 ; 
   reg __397906_397906;
   reg _397907_397907 ; 
   reg __397907_397907;
   reg _397908_397908 ; 
   reg __397908_397908;
   reg _397909_397909 ; 
   reg __397909_397909;
   reg _397910_397910 ; 
   reg __397910_397910;
   reg _397911_397911 ; 
   reg __397911_397911;
   reg _397912_397912 ; 
   reg __397912_397912;
   reg _397913_397913 ; 
   reg __397913_397913;
   reg _397914_397914 ; 
   reg __397914_397914;
   reg _397915_397915 ; 
   reg __397915_397915;
   reg _397916_397916 ; 
   reg __397916_397916;
   reg _397917_397917 ; 
   reg __397917_397917;
   reg _397918_397918 ; 
   reg __397918_397918;
   reg _397919_397919 ; 
   reg __397919_397919;
   reg _397920_397920 ; 
   reg __397920_397920;
   reg _397921_397921 ; 
   reg __397921_397921;
   reg _397922_397922 ; 
   reg __397922_397922;
   reg _397923_397923 ; 
   reg __397923_397923;
   reg _397924_397924 ; 
   reg __397924_397924;
   reg _397925_397925 ; 
   reg __397925_397925;
   reg _397926_397926 ; 
   reg __397926_397926;
   reg _397927_397927 ; 
   reg __397927_397927;
   reg _397928_397928 ; 
   reg __397928_397928;
   reg _397929_397929 ; 
   reg __397929_397929;
   reg _397930_397930 ; 
   reg __397930_397930;
   reg _397931_397931 ; 
   reg __397931_397931;
   reg _397932_397932 ; 
   reg __397932_397932;
   reg _397933_397933 ; 
   reg __397933_397933;
   reg _397934_397934 ; 
   reg __397934_397934;
   reg _397935_397935 ; 
   reg __397935_397935;
   reg _397936_397936 ; 
   reg __397936_397936;
   reg _397937_397937 ; 
   reg __397937_397937;
   reg _397938_397938 ; 
   reg __397938_397938;
   reg _397939_397939 ; 
   reg __397939_397939;
   reg _397940_397940 ; 
   reg __397940_397940;
   reg _397941_397941 ; 
   reg __397941_397941;
   reg _397942_397942 ; 
   reg __397942_397942;
   reg _397943_397943 ; 
   reg __397943_397943;
   reg _397944_397944 ; 
   reg __397944_397944;
   reg _397945_397945 ; 
   reg __397945_397945;
   reg _397946_397946 ; 
   reg __397946_397946;
   reg _397947_397947 ; 
   reg __397947_397947;
   reg _397948_397948 ; 
   reg __397948_397948;
   reg _397949_397949 ; 
   reg __397949_397949;
   reg _397950_397950 ; 
   reg __397950_397950;
   reg _397951_397951 ; 
   reg __397951_397951;
   reg _397952_397952 ; 
   reg __397952_397952;
   reg _397953_397953 ; 
   reg __397953_397953;
   reg _397954_397954 ; 
   reg __397954_397954;
   reg _397955_397955 ; 
   reg __397955_397955;
   reg _397956_397956 ; 
   reg __397956_397956;
   reg _397957_397957 ; 
   reg __397957_397957;
   reg _397958_397958 ; 
   reg __397958_397958;
   reg _397959_397959 ; 
   reg __397959_397959;
   reg _397960_397960 ; 
   reg __397960_397960;
   reg _397961_397961 ; 
   reg __397961_397961;
   reg _397962_397962 ; 
   reg __397962_397962;
   reg _397963_397963 ; 
   reg __397963_397963;
   reg _397964_397964 ; 
   reg __397964_397964;
   reg _397965_397965 ; 
   reg __397965_397965;
   reg _397966_397966 ; 
   reg __397966_397966;
   reg _397967_397967 ; 
   reg __397967_397967;
   reg _397968_397968 ; 
   reg __397968_397968;
   reg _397969_397969 ; 
   reg __397969_397969;
   reg _397970_397970 ; 
   reg __397970_397970;
   reg _397971_397971 ; 
   reg __397971_397971;
   reg _397972_397972 ; 
   reg __397972_397972;
   reg _397973_397973 ; 
   reg __397973_397973;
   reg _397974_397974 ; 
   reg __397974_397974;
   reg _397975_397975 ; 
   reg __397975_397975;
   reg _397976_397976 ; 
   reg __397976_397976;
   reg _397977_397977 ; 
   reg __397977_397977;
   reg _397978_397978 ; 
   reg __397978_397978;
   reg _397979_397979 ; 
   reg __397979_397979;
   reg _397980_397980 ; 
   reg __397980_397980;
   reg _397981_397981 ; 
   reg __397981_397981;
   reg _397982_397982 ; 
   reg __397982_397982;
   reg _397983_397983 ; 
   reg __397983_397983;
   reg _397984_397984 ; 
   reg __397984_397984;
   reg _397985_397985 ; 
   reg __397985_397985;
   reg _397986_397986 ; 
   reg __397986_397986;
   reg _397987_397987 ; 
   reg __397987_397987;
   reg _397988_397988 ; 
   reg __397988_397988;
   reg _397989_397989 ; 
   reg __397989_397989;
   reg _397990_397990 ; 
   reg __397990_397990;
   reg _397991_397991 ; 
   reg __397991_397991;
   reg _397992_397992 ; 
   reg __397992_397992;
   reg _397993_397993 ; 
   reg __397993_397993;
   reg _397994_397994 ; 
   reg __397994_397994;
   reg _397995_397995 ; 
   reg __397995_397995;
   reg _397996_397996 ; 
   reg __397996_397996;
   reg _397997_397997 ; 
   reg __397997_397997;
   reg _397998_397998 ; 
   reg __397998_397998;
   reg _397999_397999 ; 
   reg __397999_397999;
   reg _398000_398000 ; 
   reg __398000_398000;
   reg _398001_398001 ; 
   reg __398001_398001;
   reg _398002_398002 ; 
   reg __398002_398002;
   reg _398003_398003 ; 
   reg __398003_398003;
   reg _398004_398004 ; 
   reg __398004_398004;
   reg _398005_398005 ; 
   reg __398005_398005;
   reg _398006_398006 ; 
   reg __398006_398006;
   reg _398007_398007 ; 
   reg __398007_398007;
   reg _398008_398008 ; 
   reg __398008_398008;
   reg _398009_398009 ; 
   reg __398009_398009;
   reg _398010_398010 ; 
   reg __398010_398010;
   reg _398011_398011 ; 
   reg __398011_398011;
   reg _398012_398012 ; 
   reg __398012_398012;
   reg _398013_398013 ; 
   reg __398013_398013;
   reg _398014_398014 ; 
   reg __398014_398014;
   reg _398015_398015 ; 
   reg __398015_398015;
   reg _398016_398016 ; 
   reg __398016_398016;
   reg _398017_398017 ; 
   reg __398017_398017;
   reg _398018_398018 ; 
   reg __398018_398018;
   reg _398019_398019 ; 
   reg __398019_398019;
   reg _398020_398020 ; 
   reg __398020_398020;
   reg _398021_398021 ; 
   reg __398021_398021;
   reg _398022_398022 ; 
   reg __398022_398022;
   reg _398023_398023 ; 
   reg __398023_398023;
   reg _398024_398024 ; 
   reg __398024_398024;
   reg _398025_398025 ; 
   reg __398025_398025;
   reg _398026_398026 ; 
   reg __398026_398026;
   reg _398027_398027 ; 
   reg __398027_398027;
   reg _398028_398028 ; 
   reg __398028_398028;
   reg _398029_398029 ; 
   reg __398029_398029;
   reg _398030_398030 ; 
   reg __398030_398030;
   reg _398031_398031 ; 
   reg __398031_398031;
   reg _398032_398032 ; 
   reg __398032_398032;
   reg _398033_398033 ; 
   reg __398033_398033;
   reg _398034_398034 ; 
   reg __398034_398034;
   reg _398035_398035 ; 
   reg __398035_398035;
   reg _398036_398036 ; 
   reg __398036_398036;
   reg _398037_398037 ; 
   reg __398037_398037;
   reg _398038_398038 ; 
   reg __398038_398038;
   reg _398039_398039 ; 
   reg __398039_398039;
   reg _398040_398040 ; 
   reg __398040_398040;
   reg _398041_398041 ; 
   reg __398041_398041;
   reg _398042_398042 ; 
   reg __398042_398042;
   reg _398043_398043 ; 
   reg __398043_398043;
   reg _398044_398044 ; 
   reg __398044_398044;
   reg _398045_398045 ; 
   reg __398045_398045;
   reg _398046_398046 ; 
   reg __398046_398046;
   reg _398047_398047 ; 
   reg __398047_398047;
   reg _398048_398048 ; 
   reg __398048_398048;
   reg _398049_398049 ; 
   reg __398049_398049;
   reg _398050_398050 ; 
   reg __398050_398050;
   reg _398051_398051 ; 
   reg __398051_398051;
   reg _398052_398052 ; 
   reg __398052_398052;
   reg _398053_398053 ; 
   reg __398053_398053;
   reg _398054_398054 ; 
   reg __398054_398054;
   reg _398055_398055 ; 
   reg __398055_398055;
   reg _398056_398056 ; 
   reg __398056_398056;
   reg _398057_398057 ; 
   reg __398057_398057;
   reg _398058_398058 ; 
   reg __398058_398058;
   reg _398059_398059 ; 
   reg __398059_398059;
   reg _398060_398060 ; 
   reg __398060_398060;
   reg _398061_398061 ; 
   reg __398061_398061;
   reg _398062_398062 ; 
   reg __398062_398062;
   reg _398063_398063 ; 
   reg __398063_398063;
   reg _398064_398064 ; 
   reg __398064_398064;
   reg _398065_398065 ; 
   reg __398065_398065;
   reg _398066_398066 ; 
   reg __398066_398066;
   reg _398067_398067 ; 
   reg __398067_398067;
   reg _398068_398068 ; 
   reg __398068_398068;
   reg _398069_398069 ; 
   reg __398069_398069;
   reg _398070_398070 ; 
   reg __398070_398070;
   reg _398071_398071 ; 
   reg __398071_398071;
   reg _398072_398072 ; 
   reg __398072_398072;
   reg _398073_398073 ; 
   reg __398073_398073;
   reg _398074_398074 ; 
   reg __398074_398074;
   reg _398075_398075 ; 
   reg __398075_398075;
   reg _398076_398076 ; 
   reg __398076_398076;
   reg _398077_398077 ; 
   reg __398077_398077;
   reg _398078_398078 ; 
   reg __398078_398078;
   reg _398079_398079 ; 
   reg __398079_398079;
   reg _398080_398080 ; 
   reg __398080_398080;
   reg _398081_398081 ; 
   reg __398081_398081;
   reg _398082_398082 ; 
   reg __398082_398082;
   reg _398083_398083 ; 
   reg __398083_398083;
   reg _398084_398084 ; 
   reg __398084_398084;
   reg _398085_398085 ; 
   reg __398085_398085;
   reg _398086_398086 ; 
   reg __398086_398086;
   reg _398087_398087 ; 
   reg __398087_398087;
   reg _398088_398088 ; 
   reg __398088_398088;
   reg _398089_398089 ; 
   reg __398089_398089;
   reg _398090_398090 ; 
   reg __398090_398090;
   reg _398091_398091 ; 
   reg __398091_398091;
   reg _398092_398092 ; 
   reg __398092_398092;
   reg _398093_398093 ; 
   reg __398093_398093;
   reg _398094_398094 ; 
   reg __398094_398094;
   reg _398095_398095 ; 
   reg __398095_398095;
   reg _398096_398096 ; 
   reg __398096_398096;
   reg _398097_398097 ; 
   reg __398097_398097;
   reg _398098_398098 ; 
   reg __398098_398098;
   reg _398099_398099 ; 
   reg __398099_398099;
   reg _398100_398100 ; 
   reg __398100_398100;
   reg _398101_398101 ; 
   reg __398101_398101;
   reg _398102_398102 ; 
   reg __398102_398102;
   reg _398103_398103 ; 
   reg __398103_398103;
   reg _398104_398104 ; 
   reg __398104_398104;
   reg _398105_398105 ; 
   reg __398105_398105;
   reg _398106_398106 ; 
   reg __398106_398106;
   reg _398107_398107 ; 
   reg __398107_398107;
   reg _398108_398108 ; 
   reg __398108_398108;
   reg _398109_398109 ; 
   reg __398109_398109;
   reg _398110_398110 ; 
   reg __398110_398110;
   reg _398111_398111 ; 
   reg __398111_398111;
   reg _398112_398112 ; 
   reg __398112_398112;
   reg _398113_398113 ; 
   reg __398113_398113;
   reg _398114_398114 ; 
   reg __398114_398114;
   reg _398115_398115 ; 
   reg __398115_398115;
   reg _398116_398116 ; 
   reg __398116_398116;
   reg _398117_398117 ; 
   reg __398117_398117;
   reg _398118_398118 ; 
   reg __398118_398118;
   reg _398119_398119 ; 
   reg __398119_398119;
   reg _398120_398120 ; 
   reg __398120_398120;
   reg _398121_398121 ; 
   reg __398121_398121;
   reg _398122_398122 ; 
   reg __398122_398122;
   reg _398123_398123 ; 
   reg __398123_398123;
   reg _398124_398124 ; 
   reg __398124_398124;
   reg _398125_398125 ; 
   reg __398125_398125;
   reg _398126_398126 ; 
   reg __398126_398126;
   reg _398127_398127 ; 
   reg __398127_398127;
   reg _398128_398128 ; 
   reg __398128_398128;
   reg _398129_398129 ; 
   reg __398129_398129;
   reg _398130_398130 ; 
   reg __398130_398130;
   reg _398131_398131 ; 
   reg __398131_398131;
   reg _398132_398132 ; 
   reg __398132_398132;
   reg _398133_398133 ; 
   reg __398133_398133;
   reg _398134_398134 ; 
   reg __398134_398134;
   reg _398135_398135 ; 
   reg __398135_398135;
   reg _398136_398136 ; 
   reg __398136_398136;
   reg _398137_398137 ; 
   reg __398137_398137;
   reg _398138_398138 ; 
   reg __398138_398138;
   reg _398139_398139 ; 
   reg __398139_398139;
   reg _398140_398140 ; 
   reg __398140_398140;
   reg _398141_398141 ; 
   reg __398141_398141;
   reg _398142_398142 ; 
   reg __398142_398142;
   reg _398143_398143 ; 
   reg __398143_398143;
   reg _398144_398144 ; 
   reg __398144_398144;
   reg _398145_398145 ; 
   reg __398145_398145;
   reg _398146_398146 ; 
   reg __398146_398146;
   reg _398147_398147 ; 
   reg __398147_398147;
   reg _398148_398148 ; 
   reg __398148_398148;
   reg _398149_398149 ; 
   reg __398149_398149;
   reg _398150_398150 ; 
   reg __398150_398150;
   reg _398151_398151 ; 
   reg __398151_398151;
   reg _398152_398152 ; 
   reg __398152_398152;
   reg _398153_398153 ; 
   reg __398153_398153;
   reg _398154_398154 ; 
   reg __398154_398154;
   reg _398155_398155 ; 
   reg __398155_398155;
   reg _398156_398156 ; 
   reg __398156_398156;
   reg _398157_398157 ; 
   reg __398157_398157;
   reg _398158_398158 ; 
   reg __398158_398158;
   reg _398159_398159 ; 
   reg __398159_398159;
   reg _398160_398160 ; 
   reg __398160_398160;
   reg _398161_398161 ; 
   reg __398161_398161;
   reg _398162_398162 ; 
   reg __398162_398162;
   reg _398163_398163 ; 
   reg __398163_398163;
   reg _398164_398164 ; 
   reg __398164_398164;
   reg _398165_398165 ; 
   reg __398165_398165;
   reg _398166_398166 ; 
   reg __398166_398166;
   reg _398167_398167 ; 
   reg __398167_398167;
   reg _398168_398168 ; 
   reg __398168_398168;
   reg _398169_398169 ; 
   reg __398169_398169;
   reg _398170_398170 ; 
   reg __398170_398170;
   reg _398171_398171 ; 
   reg __398171_398171;
   reg _398172_398172 ; 
   reg __398172_398172;
   reg _398173_398173 ; 
   reg __398173_398173;
   reg _398174_398174 ; 
   reg __398174_398174;
   reg _398175_398175 ; 
   reg __398175_398175;
   reg _398176_398176 ; 
   reg __398176_398176;
   reg _398177_398177 ; 
   reg __398177_398177;
   reg _398178_398178 ; 
   reg __398178_398178;
   reg _398179_398179 ; 
   reg __398179_398179;
   reg _398180_398180 ; 
   reg __398180_398180;
   reg _398181_398181 ; 
   reg __398181_398181;
   reg _398182_398182 ; 
   reg __398182_398182;
   reg _398183_398183 ; 
   reg __398183_398183;
   reg _398184_398184 ; 
   reg __398184_398184;
   reg _398185_398185 ; 
   reg __398185_398185;
   reg _398186_398186 ; 
   reg __398186_398186;
   reg _398187_398187 ; 
   reg __398187_398187;
   reg _398188_398188 ; 
   reg __398188_398188;
   reg _398189_398189 ; 
   reg __398189_398189;
   reg _398190_398190 ; 
   reg __398190_398190;
   reg _398191_398191 ; 
   reg __398191_398191;
   reg _398192_398192 ; 
   reg __398192_398192;
   reg _398193_398193 ; 
   reg __398193_398193;
   reg _398194_398194 ; 
   reg __398194_398194;
   reg _398195_398195 ; 
   reg __398195_398195;
   reg _398196_398196 ; 
   reg __398196_398196;
   reg _398197_398197 ; 
   reg __398197_398197;
   reg _398198_398198 ; 
   reg __398198_398198;
   reg _398199_398199 ; 
   reg __398199_398199;
   reg _398200_398200 ; 
   reg __398200_398200;
   reg _398201_398201 ; 
   reg __398201_398201;
   reg _398202_398202 ; 
   reg __398202_398202;
   reg _398203_398203 ; 
   reg __398203_398203;
   reg _398204_398204 ; 
   reg __398204_398204;
   reg _398205_398205 ; 
   reg __398205_398205;
   reg _398206_398206 ; 
   reg __398206_398206;
   reg _398207_398207 ; 
   reg __398207_398207;
   reg _398208_398208 ; 
   reg __398208_398208;
   reg _398209_398209 ; 
   reg __398209_398209;
   reg _398210_398210 ; 
   reg __398210_398210;
   reg _398211_398211 ; 
   reg __398211_398211;
   reg _398212_398212 ; 
   reg __398212_398212;
   reg _398213_398213 ; 
   reg __398213_398213;
   reg _398214_398214 ; 
   reg __398214_398214;
   reg _398215_398215 ; 
   reg __398215_398215;
   reg _398216_398216 ; 
   reg __398216_398216;
   reg _398217_398217 ; 
   reg __398217_398217;
   reg _398218_398218 ; 
   reg __398218_398218;
   reg _398219_398219 ; 
   reg __398219_398219;
   reg _398220_398220 ; 
   reg __398220_398220;
   reg _398221_398221 ; 
   reg __398221_398221;
   reg _398222_398222 ; 
   reg __398222_398222;
   reg _398223_398223 ; 
   reg __398223_398223;
   reg _398224_398224 ; 
   reg __398224_398224;
   reg _398225_398225 ; 
   reg __398225_398225;
   reg _398226_398226 ; 
   reg __398226_398226;
   reg _398227_398227 ; 
   reg __398227_398227;
   reg _398228_398228 ; 
   reg __398228_398228;
   reg _398229_398229 ; 
   reg __398229_398229;
   reg _398230_398230 ; 
   reg __398230_398230;
   reg _398231_398231 ; 
   reg __398231_398231;
   reg _398232_398232 ; 
   reg __398232_398232;
   reg _398233_398233 ; 
   reg __398233_398233;
   reg _398234_398234 ; 
   reg __398234_398234;
   reg _398235_398235 ; 
   reg __398235_398235;
   reg _398236_398236 ; 
   reg __398236_398236;
   reg _398237_398237 ; 
   reg __398237_398237;
   reg _398238_398238 ; 
   reg __398238_398238;
   reg _398239_398239 ; 
   reg __398239_398239;
   reg _398240_398240 ; 
   reg __398240_398240;
   reg _398241_398241 ; 
   reg __398241_398241;
   reg _398242_398242 ; 
   reg __398242_398242;
   reg _398243_398243 ; 
   reg __398243_398243;
   reg _398244_398244 ; 
   reg __398244_398244;
   reg _398245_398245 ; 
   reg __398245_398245;
   reg _398246_398246 ; 
   reg __398246_398246;
   reg _398247_398247 ; 
   reg __398247_398247;
   reg _398248_398248 ; 
   reg __398248_398248;
   reg _398249_398249 ; 
   reg __398249_398249;
   reg _398250_398250 ; 
   reg __398250_398250;
   reg _398251_398251 ; 
   reg __398251_398251;
   reg _398252_398252 ; 
   reg __398252_398252;
   reg _398253_398253 ; 
   reg __398253_398253;
   reg _398254_398254 ; 
   reg __398254_398254;
   reg _398255_398255 ; 
   reg __398255_398255;
   reg _398256_398256 ; 
   reg __398256_398256;
   reg _398257_398257 ; 
   reg __398257_398257;
   reg _398258_398258 ; 
   reg __398258_398258;
   reg _398259_398259 ; 
   reg __398259_398259;
   reg _398260_398260 ; 
   reg __398260_398260;
   reg _398261_398261 ; 
   reg __398261_398261;
   reg _398262_398262 ; 
   reg __398262_398262;
   reg _398263_398263 ; 
   reg __398263_398263;
   reg _398264_398264 ; 
   reg __398264_398264;
   reg _398265_398265 ; 
   reg __398265_398265;
   reg _398266_398266 ; 
   reg __398266_398266;
   reg _398267_398267 ; 
   reg __398267_398267;
   reg _398268_398268 ; 
   reg __398268_398268;
   reg _398269_398269 ; 
   reg __398269_398269;
   reg _398270_398270 ; 
   reg __398270_398270;
   reg _398271_398271 ; 
   reg __398271_398271;
   reg _398272_398272 ; 
   reg __398272_398272;
   reg _398273_398273 ; 
   reg __398273_398273;
   reg _398274_398274 ; 
   reg __398274_398274;
   reg _398275_398275 ; 
   reg __398275_398275;
   reg _398276_398276 ; 
   reg __398276_398276;
   reg _398277_398277 ; 
   reg __398277_398277;
   reg _398278_398278 ; 
   reg __398278_398278;
   reg _398279_398279 ; 
   reg __398279_398279;
   reg _398280_398280 ; 
   reg __398280_398280;
   reg _398281_398281 ; 
   reg __398281_398281;
   reg _398282_398282 ; 
   reg __398282_398282;
   reg _398283_398283 ; 
   reg __398283_398283;
   reg _398284_398284 ; 
   reg __398284_398284;
   reg _398285_398285 ; 
   reg __398285_398285;
   reg _398286_398286 ; 
   reg __398286_398286;
   reg _398287_398287 ; 
   reg __398287_398287;
   reg _398288_398288 ; 
   reg __398288_398288;
   reg _398289_398289 ; 
   reg __398289_398289;
   reg _398290_398290 ; 
   reg __398290_398290;
   reg _398291_398291 ; 
   reg __398291_398291;
   reg _398292_398292 ; 
   reg __398292_398292;
   reg _398293_398293 ; 
   reg __398293_398293;
   reg _398294_398294 ; 
   reg __398294_398294;
   reg _398295_398295 ; 
   reg __398295_398295;
   reg _398296_398296 ; 
   reg __398296_398296;
   reg _398297_398297 ; 
   reg __398297_398297;
   reg _398298_398298 ; 
   reg __398298_398298;
   reg _398299_398299 ; 
   reg __398299_398299;
   reg _398300_398300 ; 
   reg __398300_398300;
   reg _398301_398301 ; 
   reg __398301_398301;
   reg _398302_398302 ; 
   reg __398302_398302;
   reg _398303_398303 ; 
   reg __398303_398303;
   reg _398304_398304 ; 
   reg __398304_398304;
   reg _398305_398305 ; 
   reg __398305_398305;
   reg _398306_398306 ; 
   reg __398306_398306;
   reg _398307_398307 ; 
   reg __398307_398307;
   reg _398308_398308 ; 
   reg __398308_398308;
   reg _398309_398309 ; 
   reg __398309_398309;
   reg _398310_398310 ; 
   reg __398310_398310;
   reg _398311_398311 ; 
   reg __398311_398311;
   reg _398312_398312 ; 
   reg __398312_398312;
   reg _398313_398313 ; 
   reg __398313_398313;
   reg _398314_398314 ; 
   reg __398314_398314;
   reg _398315_398315 ; 
   reg __398315_398315;
   reg _398316_398316 ; 
   reg __398316_398316;
   reg _398317_398317 ; 
   reg __398317_398317;
   reg _398318_398318 ; 
   reg __398318_398318;
   reg _398319_398319 ; 
   reg __398319_398319;
   reg _398320_398320 ; 
   reg __398320_398320;
   reg _398321_398321 ; 
   reg __398321_398321;
   reg _398322_398322 ; 
   reg __398322_398322;
   reg _398323_398323 ; 
   reg __398323_398323;
   reg _398324_398324 ; 
   reg __398324_398324;
   reg _398325_398325 ; 
   reg __398325_398325;
   reg _398326_398326 ; 
   reg __398326_398326;
   reg _398327_398327 ; 
   reg __398327_398327;
   reg _398328_398328 ; 
   reg __398328_398328;
   reg _398329_398329 ; 
   reg __398329_398329;
   reg _398330_398330 ; 
   reg __398330_398330;
   reg _398331_398331 ; 
   reg __398331_398331;
   reg _398332_398332 ; 
   reg __398332_398332;
   reg _398333_398333 ; 
   reg __398333_398333;
   reg _398334_398334 ; 
   reg __398334_398334;
   reg _398335_398335 ; 
   reg __398335_398335;
   reg _398336_398336 ; 
   reg __398336_398336;
   reg _398337_398337 ; 
   reg __398337_398337;
   reg _398338_398338 ; 
   reg __398338_398338;
   reg _398339_398339 ; 
   reg __398339_398339;
   reg _398340_398340 ; 
   reg __398340_398340;
   reg _398341_398341 ; 
   reg __398341_398341;
   reg _398342_398342 ; 
   reg __398342_398342;
   reg _398343_398343 ; 
   reg __398343_398343;
   reg _398344_398344 ; 
   reg __398344_398344;
   reg _398345_398345 ; 
   reg __398345_398345;
   reg _398346_398346 ; 
   reg __398346_398346;
   reg _398347_398347 ; 
   reg __398347_398347;
   reg _398348_398348 ; 
   reg __398348_398348;
   reg _398349_398349 ; 
   reg __398349_398349;
   reg _398350_398350 ; 
   reg __398350_398350;
   reg _398351_398351 ; 
   reg __398351_398351;
   reg _398352_398352 ; 
   reg __398352_398352;
   reg _398353_398353 ; 
   reg __398353_398353;
   reg _398354_398354 ; 
   reg __398354_398354;
   reg _398355_398355 ; 
   reg __398355_398355;
   reg _398356_398356 ; 
   reg __398356_398356;
   reg _398357_398357 ; 
   reg __398357_398357;
   reg _398358_398358 ; 
   reg __398358_398358;
   reg _398359_398359 ; 
   reg __398359_398359;
   reg _398360_398360 ; 
   reg __398360_398360;
   reg _398361_398361 ; 
   reg __398361_398361;
   reg _398362_398362 ; 
   reg __398362_398362;
   reg _398363_398363 ; 
   reg __398363_398363;
   reg _398364_398364 ; 
   reg __398364_398364;
   reg _398365_398365 ; 
   reg __398365_398365;
   reg _398366_398366 ; 
   reg __398366_398366;
   reg _398367_398367 ; 
   reg __398367_398367;
   reg _398368_398368 ; 
   reg __398368_398368;
   reg _398369_398369 ; 
   reg __398369_398369;
   reg _398370_398370 ; 
   reg __398370_398370;
   reg _398371_398371 ; 
   reg __398371_398371;
   reg _398372_398372 ; 
   reg __398372_398372;
   reg _398373_398373 ; 
   reg __398373_398373;
   reg _398374_398374 ; 
   reg __398374_398374;
   reg _398375_398375 ; 
   reg __398375_398375;
   reg _398376_398376 ; 
   reg __398376_398376;
   reg _398377_398377 ; 
   reg __398377_398377;
   reg _398378_398378 ; 
   reg __398378_398378;
   reg _398379_398379 ; 
   reg __398379_398379;
   reg _398380_398380 ; 
   reg __398380_398380;
   reg _398381_398381 ; 
   reg __398381_398381;
   reg _398382_398382 ; 
   reg __398382_398382;
   reg _398383_398383 ; 
   reg __398383_398383;
   reg _398384_398384 ; 
   reg __398384_398384;
   reg _398385_398385 ; 
   reg __398385_398385;
   reg _398386_398386 ; 
   reg __398386_398386;
   reg _398387_398387 ; 
   reg __398387_398387;
   reg _398388_398388 ; 
   reg __398388_398388;
   reg _398389_398389 ; 
   reg __398389_398389;
   reg _398390_398390 ; 
   reg __398390_398390;
   reg _398391_398391 ; 
   reg __398391_398391;
   reg _398392_398392 ; 
   reg __398392_398392;
   reg _398393_398393 ; 
   reg __398393_398393;
   reg _398394_398394 ; 
   reg __398394_398394;
   reg _398395_398395 ; 
   reg __398395_398395;
   reg _398396_398396 ; 
   reg __398396_398396;
   reg _398397_398397 ; 
   reg __398397_398397;
   reg _398398_398398 ; 
   reg __398398_398398;
   reg _398399_398399 ; 
   reg __398399_398399;
   reg _398400_398400 ; 
   reg __398400_398400;
   reg _398401_398401 ; 
   reg __398401_398401;
   reg _398402_398402 ; 
   reg __398402_398402;
   reg _398403_398403 ; 
   reg __398403_398403;
   reg _398404_398404 ; 
   reg __398404_398404;
   reg _398405_398405 ; 
   reg __398405_398405;
   reg _398406_398406 ; 
   reg __398406_398406;
   reg _398407_398407 ; 
   reg __398407_398407;
   reg _398408_398408 ; 
   reg __398408_398408;
   reg _398409_398409 ; 
   reg __398409_398409;
   reg _398410_398410 ; 
   reg __398410_398410;
   reg _398411_398411 ; 
   reg __398411_398411;
   reg _398412_398412 ; 
   reg __398412_398412;
   reg _398413_398413 ; 
   reg __398413_398413;
   reg _398414_398414 ; 
   reg __398414_398414;
   reg _398415_398415 ; 
   reg __398415_398415;
   reg _398416_398416 ; 
   reg __398416_398416;
   reg _398417_398417 ; 
   reg __398417_398417;
   reg _398418_398418 ; 
   reg __398418_398418;
   reg _398419_398419 ; 
   reg __398419_398419;
   reg _398420_398420 ; 
   reg __398420_398420;
   reg _398421_398421 ; 
   reg __398421_398421;
   reg _398422_398422 ; 
   reg __398422_398422;
   reg _398423_398423 ; 
   reg __398423_398423;
   reg _398424_398424 ; 
   reg __398424_398424;
   reg _398425_398425 ; 
   reg __398425_398425;
   reg _398426_398426 ; 
   reg __398426_398426;
   reg _398427_398427 ; 
   reg __398427_398427;
   reg _398428_398428 ; 
   reg __398428_398428;
   reg _398429_398429 ; 
   reg __398429_398429;
   reg _398430_398430 ; 
   reg __398430_398430;
   reg _398431_398431 ; 
   reg __398431_398431;
   reg _398432_398432 ; 
   reg __398432_398432;
   reg _398433_398433 ; 
   reg __398433_398433;
   reg _398434_398434 ; 
   reg __398434_398434;
   reg _398435_398435 ; 
   reg __398435_398435;
   reg _398436_398436 ; 
   reg __398436_398436;
   reg _398437_398437 ; 
   reg __398437_398437;
   reg _398438_398438 ; 
   reg __398438_398438;
   reg _398439_398439 ; 
   reg __398439_398439;
   reg _398440_398440 ; 
   reg __398440_398440;
   reg _398441_398441 ; 
   reg __398441_398441;
   reg _398442_398442 ; 
   reg __398442_398442;
   reg _398443_398443 ; 
   reg __398443_398443;
   reg _398444_398444 ; 
   reg __398444_398444;
   reg _398445_398445 ; 
   reg __398445_398445;
   reg _398446_398446 ; 
   reg __398446_398446;
   reg _398447_398447 ; 
   reg __398447_398447;
   reg _398448_398448 ; 
   reg __398448_398448;
   reg _398449_398449 ; 
   reg __398449_398449;
   reg _398450_398450 ; 
   reg __398450_398450;
   reg _398451_398451 ; 
   reg __398451_398451;
   reg _398452_398452 ; 
   reg __398452_398452;
   reg _398453_398453 ; 
   reg __398453_398453;
   reg _398454_398454 ; 
   reg __398454_398454;
   reg _398455_398455 ; 
   reg __398455_398455;
   reg _398456_398456 ; 
   reg __398456_398456;
   reg _398457_398457 ; 
   reg __398457_398457;
   reg _398458_398458 ; 
   reg __398458_398458;
   reg _398459_398459 ; 
   reg __398459_398459;
   reg _398460_398460 ; 
   reg __398460_398460;
   reg _398461_398461 ; 
   reg __398461_398461;
   reg _398462_398462 ; 
   reg __398462_398462;
   reg _398463_398463 ; 
   reg __398463_398463;
   reg _398464_398464 ; 
   reg __398464_398464;
   reg _398465_398465 ; 
   reg __398465_398465;
   reg _398466_398466 ; 
   reg __398466_398466;
   reg _398467_398467 ; 
   reg __398467_398467;
   reg _398468_398468 ; 
   reg __398468_398468;
   reg _398469_398469 ; 
   reg __398469_398469;
   reg _398470_398470 ; 
   reg __398470_398470;
   reg _398471_398471 ; 
   reg __398471_398471;
   reg _398472_398472 ; 
   reg __398472_398472;
   reg _398473_398473 ; 
   reg __398473_398473;
   reg _398474_398474 ; 
   reg __398474_398474;
   reg _398475_398475 ; 
   reg __398475_398475;
   reg _398476_398476 ; 
   reg __398476_398476;
   reg _398477_398477 ; 
   reg __398477_398477;
   reg _398478_398478 ; 
   reg __398478_398478;
   reg _398479_398479 ; 
   reg __398479_398479;
   reg _398480_398480 ; 
   reg __398480_398480;
   reg _398481_398481 ; 
   reg __398481_398481;
   reg _398482_398482 ; 
   reg __398482_398482;
   reg _398483_398483 ; 
   reg __398483_398483;
   reg _398484_398484 ; 
   reg __398484_398484;
   reg _398485_398485 ; 
   reg __398485_398485;
   reg _398486_398486 ; 
   reg __398486_398486;
   reg _398487_398487 ; 
   reg __398487_398487;
   reg _398488_398488 ; 
   reg __398488_398488;
   reg _398489_398489 ; 
   reg __398489_398489;
   reg _398490_398490 ; 
   reg __398490_398490;
   reg _398491_398491 ; 
   reg __398491_398491;
   reg _398492_398492 ; 
   reg __398492_398492;
   reg _398493_398493 ; 
   reg __398493_398493;
   reg _398494_398494 ; 
   reg __398494_398494;
   reg _398495_398495 ; 
   reg __398495_398495;
   reg _398496_398496 ; 
   reg __398496_398496;
   reg _398497_398497 ; 
   reg __398497_398497;
   reg _398498_398498 ; 
   reg __398498_398498;
   reg _398499_398499 ; 
   reg __398499_398499;
   reg _398500_398500 ; 
   reg __398500_398500;
   reg _398501_398501 ; 
   reg __398501_398501;
   reg _398502_398502 ; 
   reg __398502_398502;
   reg _398503_398503 ; 
   reg __398503_398503;
   reg _398504_398504 ; 
   reg __398504_398504;
   reg _398505_398505 ; 
   reg __398505_398505;
   reg _398506_398506 ; 
   reg __398506_398506;
   reg _398507_398507 ; 
   reg __398507_398507;
   reg _398508_398508 ; 
   reg __398508_398508;
   reg _398509_398509 ; 
   reg __398509_398509;
   reg _398510_398510 ; 
   reg __398510_398510;
   reg _398511_398511 ; 
   reg __398511_398511;
   reg _398512_398512 ; 
   reg __398512_398512;
   reg _398513_398513 ; 
   reg __398513_398513;
   reg _398514_398514 ; 
   reg __398514_398514;
   reg _398515_398515 ; 
   reg __398515_398515;
   reg _398516_398516 ; 
   reg __398516_398516;
   reg _398517_398517 ; 
   reg __398517_398517;
   reg _398518_398518 ; 
   reg __398518_398518;
   reg _398519_398519 ; 
   reg __398519_398519;
   reg _398520_398520 ; 
   reg __398520_398520;
   reg _398521_398521 ; 
   reg __398521_398521;
   reg _398522_398522 ; 
   reg __398522_398522;
   reg _398523_398523 ; 
   reg __398523_398523;
   reg _398524_398524 ; 
   reg __398524_398524;
   reg _398525_398525 ; 
   reg __398525_398525;
   reg _398526_398526 ; 
   reg __398526_398526;
   reg _398527_398527 ; 
   reg __398527_398527;
   reg _398528_398528 ; 
   reg __398528_398528;
   reg _398529_398529 ; 
   reg __398529_398529;
   reg _398530_398530 ; 
   reg __398530_398530;
   reg _398531_398531 ; 
   reg __398531_398531;
   reg _398532_398532 ; 
   reg __398532_398532;
   reg _398533_398533 ; 
   reg __398533_398533;
   reg _398534_398534 ; 
   reg __398534_398534;
   reg _398535_398535 ; 
   reg __398535_398535;
   reg _398536_398536 ; 
   reg __398536_398536;
   reg _398537_398537 ; 
   reg __398537_398537;
   reg _398538_398538 ; 
   reg __398538_398538;
   reg _398539_398539 ; 
   reg __398539_398539;
   reg _398540_398540 ; 
   reg __398540_398540;
   reg _398541_398541 ; 
   reg __398541_398541;
   reg _398542_398542 ; 
   reg __398542_398542;
   reg _398543_398543 ; 
   reg __398543_398543;
   reg _398544_398544 ; 
   reg __398544_398544;
   reg _398545_398545 ; 
   reg __398545_398545;
   reg _398546_398546 ; 
   reg __398546_398546;
   reg _398547_398547 ; 
   reg __398547_398547;
   reg _398548_398548 ; 
   reg __398548_398548;
   reg _398549_398549 ; 
   reg __398549_398549;
   reg _398550_398550 ; 
   reg __398550_398550;
   reg _398551_398551 ; 
   reg __398551_398551;
   reg _398552_398552 ; 
   reg __398552_398552;
   reg _398553_398553 ; 
   reg __398553_398553;
   reg _398554_398554 ; 
   reg __398554_398554;
   reg _398555_398555 ; 
   reg __398555_398555;
   reg _398556_398556 ; 
   reg __398556_398556;
   reg _398557_398557 ; 
   reg __398557_398557;
   reg _398558_398558 ; 
   reg __398558_398558;
   reg _398559_398559 ; 
   reg __398559_398559;
   reg _398560_398560 ; 
   reg __398560_398560;
   reg _398561_398561 ; 
   reg __398561_398561;
   reg _398562_398562 ; 
   reg __398562_398562;
   reg _398563_398563 ; 
   reg __398563_398563;
   reg _398564_398564 ; 
   reg __398564_398564;
   reg _398565_398565 ; 
   reg __398565_398565;
   reg _398566_398566 ; 
   reg __398566_398566;
   reg _398567_398567 ; 
   reg __398567_398567;
   reg _398568_398568 ; 
   reg __398568_398568;
   reg _398569_398569 ; 
   reg __398569_398569;
   reg _398570_398570 ; 
   reg __398570_398570;
   reg _398571_398571 ; 
   reg __398571_398571;
   reg _398572_398572 ; 
   reg __398572_398572;
   reg _398573_398573 ; 
   reg __398573_398573;
   reg _398574_398574 ; 
   reg __398574_398574;
   reg _398575_398575 ; 
   reg __398575_398575;
   reg _398576_398576 ; 
   reg __398576_398576;
   reg _398577_398577 ; 
   reg __398577_398577;
   reg _398578_398578 ; 
   reg __398578_398578;
   reg _398579_398579 ; 
   reg __398579_398579;
   reg _398580_398580 ; 
   reg __398580_398580;
   reg _398581_398581 ; 
   reg __398581_398581;
   reg _398582_398582 ; 
   reg __398582_398582;
   reg _398583_398583 ; 
   reg __398583_398583;
   reg _398584_398584 ; 
   reg __398584_398584;
   reg _398585_398585 ; 
   reg __398585_398585;
   reg _398586_398586 ; 
   reg __398586_398586;
   reg _398587_398587 ; 
   reg __398587_398587;
   reg _398588_398588 ; 
   reg __398588_398588;
   reg _398589_398589 ; 
   reg __398589_398589;
   reg _398590_398590 ; 
   reg __398590_398590;
   reg _398591_398591 ; 
   reg __398591_398591;
   reg _398592_398592 ; 
   reg __398592_398592;
   reg _398593_398593 ; 
   reg __398593_398593;
   reg _398594_398594 ; 
   reg __398594_398594;
   reg _398595_398595 ; 
   reg __398595_398595;
   reg _398596_398596 ; 
   reg __398596_398596;
   reg _398597_398597 ; 
   reg __398597_398597;
   reg _398598_398598 ; 
   reg __398598_398598;
   reg _398599_398599 ; 
   reg __398599_398599;
   reg _398600_398600 ; 
   reg __398600_398600;
   reg _398601_398601 ; 
   reg __398601_398601;
   reg _398602_398602 ; 
   reg __398602_398602;
   reg _398603_398603 ; 
   reg __398603_398603;
   reg _398604_398604 ; 
   reg __398604_398604;
   reg _398605_398605 ; 
   reg __398605_398605;
   reg _398606_398606 ; 
   reg __398606_398606;
   reg _398607_398607 ; 
   reg __398607_398607;
   reg _398608_398608 ; 
   reg __398608_398608;
   reg _398609_398609 ; 
   reg __398609_398609;
   reg _398610_398610 ; 
   reg __398610_398610;
   reg _398611_398611 ; 
   reg __398611_398611;
   reg _398612_398612 ; 
   reg __398612_398612;
   reg _398613_398613 ; 
   reg __398613_398613;
   reg _398614_398614 ; 
   reg __398614_398614;
   reg _398615_398615 ; 
   reg __398615_398615;
   reg _398616_398616 ; 
   reg __398616_398616;
   reg _398617_398617 ; 
   reg __398617_398617;
   reg _398618_398618 ; 
   reg __398618_398618;
   reg _398619_398619 ; 
   reg __398619_398619;
   reg _398620_398620 ; 
   reg __398620_398620;
   reg _398621_398621 ; 
   reg __398621_398621;
   reg _398622_398622 ; 
   reg __398622_398622;
   reg _398623_398623 ; 
   reg __398623_398623;
   reg _398624_398624 ; 
   reg __398624_398624;
   reg _398625_398625 ; 
   reg __398625_398625;
   reg _398626_398626 ; 
   reg __398626_398626;
   reg _398627_398627 ; 
   reg __398627_398627;
   reg _398628_398628 ; 
   reg __398628_398628;
   reg _398629_398629 ; 
   reg __398629_398629;
   reg _398630_398630 ; 
   reg __398630_398630;
   reg _398631_398631 ; 
   reg __398631_398631;
   reg _398632_398632 ; 
   reg __398632_398632;
   reg _398633_398633 ; 
   reg __398633_398633;
   reg _398634_398634 ; 
   reg __398634_398634;
   reg _398635_398635 ; 
   reg __398635_398635;
   reg _398636_398636 ; 
   reg __398636_398636;
   reg _398637_398637 ; 
   reg __398637_398637;
   reg _398638_398638 ; 
   reg __398638_398638;
   reg _398639_398639 ; 
   reg __398639_398639;
   reg _398640_398640 ; 
   reg __398640_398640;
   reg _398641_398641 ; 
   reg __398641_398641;
   reg _398642_398642 ; 
   reg __398642_398642;
   reg _398643_398643 ; 
   reg __398643_398643;
   reg _398644_398644 ; 
   reg __398644_398644;
   reg _398645_398645 ; 
   reg __398645_398645;
   reg _398646_398646 ; 
   reg __398646_398646;
   reg _398647_398647 ; 
   reg __398647_398647;
   reg _398648_398648 ; 
   reg __398648_398648;
   reg _398649_398649 ; 
   reg __398649_398649;
   reg _398650_398650 ; 
   reg __398650_398650;
   reg _398651_398651 ; 
   reg __398651_398651;
   reg _398652_398652 ; 
   reg __398652_398652;
   reg _398653_398653 ; 
   reg __398653_398653;
   reg _398654_398654 ; 
   reg __398654_398654;
   reg _398655_398655 ; 
   reg __398655_398655;
   reg _398656_398656 ; 
   reg __398656_398656;
   reg _398657_398657 ; 
   reg __398657_398657;
   reg _398658_398658 ; 
   reg __398658_398658;
   reg _398659_398659 ; 
   reg __398659_398659;
   reg _398660_398660 ; 
   reg __398660_398660;
   reg _398661_398661 ; 
   reg __398661_398661;
   reg _398662_398662 ; 
   reg __398662_398662;
   reg _398663_398663 ; 
   reg __398663_398663;
   reg _398664_398664 ; 
   reg __398664_398664;
   reg _398665_398665 ; 
   reg __398665_398665;
   reg _398666_398666 ; 
   reg __398666_398666;
   reg _398667_398667 ; 
   reg __398667_398667;
   reg _398668_398668 ; 
   reg __398668_398668;
   reg _398669_398669 ; 
   reg __398669_398669;
   reg _398670_398670 ; 
   reg __398670_398670;
   reg _398671_398671 ; 
   reg __398671_398671;
   reg _398672_398672 ; 
   reg __398672_398672;
   reg _398673_398673 ; 
   reg __398673_398673;
   reg _398674_398674 ; 
   reg __398674_398674;
   reg _398675_398675 ; 
   reg __398675_398675;
   reg _398676_398676 ; 
   reg __398676_398676;
   reg _398677_398677 ; 
   reg __398677_398677;
   reg _398678_398678 ; 
   reg __398678_398678;
   reg _398679_398679 ; 
   reg __398679_398679;
   reg _398680_398680 ; 
   reg __398680_398680;
   reg _398681_398681 ; 
   reg __398681_398681;
   reg _398682_398682 ; 
   reg __398682_398682;
   reg _398683_398683 ; 
   reg __398683_398683;
   reg _398684_398684 ; 
   reg __398684_398684;
   reg _398685_398685 ; 
   reg __398685_398685;
   reg _398686_398686 ; 
   reg __398686_398686;
   reg _398687_398687 ; 
   reg __398687_398687;
   reg _398688_398688 ; 
   reg __398688_398688;
   reg _398689_398689 ; 
   reg __398689_398689;
   reg _398690_398690 ; 
   reg __398690_398690;
   reg _398691_398691 ; 
   reg __398691_398691;
   reg _398692_398692 ; 
   reg __398692_398692;
   reg _398693_398693 ; 
   reg __398693_398693;
   reg _398694_398694 ; 
   reg __398694_398694;
   reg _398695_398695 ; 
   reg __398695_398695;
   reg _398696_398696 ; 
   reg __398696_398696;
   reg _398697_398697 ; 
   reg __398697_398697;
   reg _398698_398698 ; 
   reg __398698_398698;
   reg _398699_398699 ; 
   reg __398699_398699;
   reg _398700_398700 ; 
   reg __398700_398700;
   reg _398701_398701 ; 
   reg __398701_398701;
   reg _398702_398702 ; 
   reg __398702_398702;
   reg _398703_398703 ; 
   reg __398703_398703;
   reg _398704_398704 ; 
   reg __398704_398704;
   reg _398705_398705 ; 
   reg __398705_398705;
   reg _398706_398706 ; 
   reg __398706_398706;
   reg _398707_398707 ; 
   reg __398707_398707;
   reg _398708_398708 ; 
   reg __398708_398708;
   reg _398709_398709 ; 
   reg __398709_398709;
   reg _398710_398710 ; 
   reg __398710_398710;
   reg _398711_398711 ; 
   reg __398711_398711;
   reg _398712_398712 ; 
   reg __398712_398712;
   reg _398713_398713 ; 
   reg __398713_398713;
   reg _398714_398714 ; 
   reg __398714_398714;
   reg _398715_398715 ; 
   reg __398715_398715;
   reg _398716_398716 ; 
   reg __398716_398716;
   reg _398717_398717 ; 
   reg __398717_398717;
   reg _398718_398718 ; 
   reg __398718_398718;
   reg _398719_398719 ; 
   reg __398719_398719;
   reg _398720_398720 ; 
   reg __398720_398720;
   reg _398721_398721 ; 
   reg __398721_398721;
   reg _398722_398722 ; 
   reg __398722_398722;
   reg _398723_398723 ; 
   reg __398723_398723;
   reg _398724_398724 ; 
   reg __398724_398724;
   reg _398725_398725 ; 
   reg __398725_398725;
   reg _398726_398726 ; 
   reg __398726_398726;
   reg _398727_398727 ; 
   reg __398727_398727;
   reg _398728_398728 ; 
   reg __398728_398728;
   reg _398729_398729 ; 
   reg __398729_398729;
   reg _398730_398730 ; 
   reg __398730_398730;
   reg _398731_398731 ; 
   reg __398731_398731;
   reg _398732_398732 ; 
   reg __398732_398732;
   reg _398733_398733 ; 
   reg __398733_398733;
   reg _398734_398734 ; 
   reg __398734_398734;
   reg _398735_398735 ; 
   reg __398735_398735;
   reg _398736_398736 ; 
   reg __398736_398736;
   reg _398737_398737 ; 
   reg __398737_398737;
   reg _398738_398738 ; 
   reg __398738_398738;
   reg _398739_398739 ; 
   reg __398739_398739;
   reg _398740_398740 ; 
   reg __398740_398740;
   reg _398741_398741 ; 
   reg __398741_398741;
   reg _398742_398742 ; 
   reg __398742_398742;
   reg _398743_398743 ; 
   reg __398743_398743;
   reg _398744_398744 ; 
   reg __398744_398744;
   reg _398745_398745 ; 
   reg __398745_398745;
   reg _398746_398746 ; 
   reg __398746_398746;
   reg _398747_398747 ; 
   reg __398747_398747;
   reg _398748_398748 ; 
   reg __398748_398748;
   reg _398749_398749 ; 
   reg __398749_398749;
   reg _398750_398750 ; 
   reg __398750_398750;
   reg _398751_398751 ; 
   reg __398751_398751;
   reg _398752_398752 ; 
   reg __398752_398752;
   reg _398753_398753 ; 
   reg __398753_398753;
   reg _398754_398754 ; 
   reg __398754_398754;
   reg _398755_398755 ; 
   reg __398755_398755;
   reg _398756_398756 ; 
   reg __398756_398756;
   reg _398757_398757 ; 
   reg __398757_398757;
   reg _398758_398758 ; 
   reg __398758_398758;
   reg _398759_398759 ; 
   reg __398759_398759;
   reg _398760_398760 ; 
   reg __398760_398760;
   reg _398761_398761 ; 
   reg __398761_398761;
   reg _398762_398762 ; 
   reg __398762_398762;
   reg _398763_398763 ; 
   reg __398763_398763;
   reg _398764_398764 ; 
   reg __398764_398764;
   reg _398765_398765 ; 
   reg __398765_398765;
   reg _398766_398766 ; 
   reg __398766_398766;
   reg _398767_398767 ; 
   reg __398767_398767;
   reg _398768_398768 ; 
   reg __398768_398768;
   reg _398769_398769 ; 
   reg __398769_398769;
   reg _398770_398770 ; 
   reg __398770_398770;
   reg _398771_398771 ; 
   reg __398771_398771;
   reg _398772_398772 ; 
   reg __398772_398772;
   reg _398773_398773 ; 
   reg __398773_398773;
   reg _398774_398774 ; 
   reg __398774_398774;
   reg _398775_398775 ; 
   reg __398775_398775;
   reg _398776_398776 ; 
   reg __398776_398776;
   reg _398777_398777 ; 
   reg __398777_398777;
   reg _398778_398778 ; 
   reg __398778_398778;
   reg _398779_398779 ; 
   reg __398779_398779;
   reg _398780_398780 ; 
   reg __398780_398780;
   reg _398781_398781 ; 
   reg __398781_398781;
   reg _398782_398782 ; 
   reg __398782_398782;
   reg _398783_398783 ; 
   reg __398783_398783;
   reg _398784_398784 ; 
   reg __398784_398784;
   reg _398785_398785 ; 
   reg __398785_398785;
   reg _398786_398786 ; 
   reg __398786_398786;
   reg _398787_398787 ; 
   reg __398787_398787;
   reg _398788_398788 ; 
   reg __398788_398788;
   reg _398789_398789 ; 
   reg __398789_398789;
   reg _398790_398790 ; 
   reg __398790_398790;
   reg _398791_398791 ; 
   reg __398791_398791;
   reg _398792_398792 ; 
   reg __398792_398792;
   reg _398793_398793 ; 
   reg __398793_398793;
   reg _398794_398794 ; 
   reg __398794_398794;
   reg _398795_398795 ; 
   reg __398795_398795;
   reg _398796_398796 ; 
   reg __398796_398796;
   reg _398797_398797 ; 
   reg __398797_398797;
   reg _398798_398798 ; 
   reg __398798_398798;
   reg _398799_398799 ; 
   reg __398799_398799;
   reg _398800_398800 ; 
   reg __398800_398800;
   reg _398801_398801 ; 
   reg __398801_398801;
   reg _398802_398802 ; 
   reg __398802_398802;
   reg _398803_398803 ; 
   reg __398803_398803;
   reg _398804_398804 ; 
   reg __398804_398804;
   reg _398805_398805 ; 
   reg __398805_398805;
   reg _398806_398806 ; 
   reg __398806_398806;
   reg _398807_398807 ; 
   reg __398807_398807;
   reg _398808_398808 ; 
   reg __398808_398808;
   reg _398809_398809 ; 
   reg __398809_398809;
   reg _398810_398810 ; 
   reg __398810_398810;
   reg _398811_398811 ; 
   reg __398811_398811;
   reg _398812_398812 ; 
   reg __398812_398812;
   reg _398813_398813 ; 
   reg __398813_398813;
   reg _398814_398814 ; 
   reg __398814_398814;
   reg _398815_398815 ; 
   reg __398815_398815;
   reg _398816_398816 ; 
   reg __398816_398816;
   reg _398817_398817 ; 
   reg __398817_398817;
   reg _398818_398818 ; 
   reg __398818_398818;
   reg _398819_398819 ; 
   reg __398819_398819;
   reg _398820_398820 ; 
   reg __398820_398820;
   reg _398821_398821 ; 
   reg __398821_398821;
   reg _398822_398822 ; 
   reg __398822_398822;
   reg _398823_398823 ; 
   reg __398823_398823;
   reg _398824_398824 ; 
   reg __398824_398824;
   reg _398825_398825 ; 
   reg __398825_398825;
   reg _398826_398826 ; 
   reg __398826_398826;
   reg _398827_398827 ; 
   reg __398827_398827;
   reg _398828_398828 ; 
   reg __398828_398828;
   reg _398829_398829 ; 
   reg __398829_398829;
   reg _398830_398830 ; 
   reg __398830_398830;
   reg _398831_398831 ; 
   reg __398831_398831;
   reg _398832_398832 ; 
   reg __398832_398832;
   reg _398833_398833 ; 
   reg __398833_398833;
   reg _398834_398834 ; 
   reg __398834_398834;
   reg _398835_398835 ; 
   reg __398835_398835;
   reg _398836_398836 ; 
   reg __398836_398836;
   reg _398837_398837 ; 
   reg __398837_398837;
   reg _398838_398838 ; 
   reg __398838_398838;
   reg _398839_398839 ; 
   reg __398839_398839;
   reg _398840_398840 ; 
   reg __398840_398840;
   reg _398841_398841 ; 
   reg __398841_398841;
   reg _398842_398842 ; 
   reg __398842_398842;
   reg _398843_398843 ; 
   reg __398843_398843;
   reg _398844_398844 ; 
   reg __398844_398844;
   reg _398845_398845 ; 
   reg __398845_398845;
   reg _398846_398846 ; 
   reg __398846_398846;
   reg _398847_398847 ; 
   reg __398847_398847;
   reg _398848_398848 ; 
   reg __398848_398848;
   reg _398849_398849 ; 
   reg __398849_398849;
   reg _398850_398850 ; 
   reg __398850_398850;
   reg _398851_398851 ; 
   reg __398851_398851;
   reg _398852_398852 ; 
   reg __398852_398852;
   reg _398853_398853 ; 
   reg __398853_398853;
   reg _398854_398854 ; 
   reg __398854_398854;
   reg _398855_398855 ; 
   reg __398855_398855;
   reg _398856_398856 ; 
   reg __398856_398856;
   reg _398857_398857 ; 
   reg __398857_398857;
   reg _398858_398858 ; 
   reg __398858_398858;
   reg _398859_398859 ; 
   reg __398859_398859;
   reg _398860_398860 ; 
   reg __398860_398860;
   reg _398861_398861 ; 
   reg __398861_398861;
   reg _398862_398862 ; 
   reg __398862_398862;
   reg _398863_398863 ; 
   reg __398863_398863;
   reg _398864_398864 ; 
   reg __398864_398864;
   reg _398865_398865 ; 
   reg __398865_398865;
   reg _398866_398866 ; 
   reg __398866_398866;
   reg _398867_398867 ; 
   reg __398867_398867;
   reg _398868_398868 ; 
   reg __398868_398868;
   reg _398869_398869 ; 
   reg __398869_398869;
   reg _398870_398870 ; 
   reg __398870_398870;
   reg _398871_398871 ; 
   reg __398871_398871;
   reg _398872_398872 ; 
   reg __398872_398872;
   reg _398873_398873 ; 
   reg __398873_398873;
   reg _398874_398874 ; 
   reg __398874_398874;
   reg _398875_398875 ; 
   reg __398875_398875;
   reg _398876_398876 ; 
   reg __398876_398876;
   reg _398877_398877 ; 
   reg __398877_398877;
   reg _398878_398878 ; 
   reg __398878_398878;
   reg _398879_398879 ; 
   reg __398879_398879;
   reg _398880_398880 ; 
   reg __398880_398880;
   reg _398881_398881 ; 
   reg __398881_398881;
   reg _398882_398882 ; 
   reg __398882_398882;
   reg _398883_398883 ; 
   reg __398883_398883;
   reg _398884_398884 ; 
   reg __398884_398884;
   reg _398885_398885 ; 
   reg __398885_398885;
   reg _398886_398886 ; 
   reg __398886_398886;
   reg _398887_398887 ; 
   reg __398887_398887;
   reg _398888_398888 ; 
   reg __398888_398888;
   reg _398889_398889 ; 
   reg __398889_398889;
   reg _398890_398890 ; 
   reg __398890_398890;
   reg _398891_398891 ; 
   reg __398891_398891;
   reg _398892_398892 ; 
   reg __398892_398892;
   reg _398893_398893 ; 
   reg __398893_398893;
   reg _398894_398894 ; 
   reg __398894_398894;
   reg _398895_398895 ; 
   reg __398895_398895;
   reg _398896_398896 ; 
   reg __398896_398896;
   reg _398897_398897 ; 
   reg __398897_398897;
   reg _398898_398898 ; 
   reg __398898_398898;
   reg _398899_398899 ; 
   reg __398899_398899;
   reg _398900_398900 ; 
   reg __398900_398900;
   reg _398901_398901 ; 
   reg __398901_398901;
   reg _398902_398902 ; 
   reg __398902_398902;
   reg _398903_398903 ; 
   reg __398903_398903;
   reg _398904_398904 ; 
   reg __398904_398904;
   reg _398905_398905 ; 
   reg __398905_398905;
   reg _398906_398906 ; 
   reg __398906_398906;
   reg _398907_398907 ; 
   reg __398907_398907;
   reg _398908_398908 ; 
   reg __398908_398908;
   reg _398909_398909 ; 
   reg __398909_398909;
   reg _398910_398910 ; 
   reg __398910_398910;
   reg _398911_398911 ; 
   reg __398911_398911;
   reg _398912_398912 ; 
   reg __398912_398912;
   reg _398913_398913 ; 
   reg __398913_398913;
   reg _398914_398914 ; 
   reg __398914_398914;
   reg _398915_398915 ; 
   reg __398915_398915;
   reg _398916_398916 ; 
   reg __398916_398916;
   reg _398917_398917 ; 
   reg __398917_398917;
   reg _398918_398918 ; 
   reg __398918_398918;
   reg _398919_398919 ; 
   reg __398919_398919;
   reg _398920_398920 ; 
   reg __398920_398920;
   reg _398921_398921 ; 
   reg __398921_398921;
   reg _398922_398922 ; 
   reg __398922_398922;
   reg _398923_398923 ; 
   reg __398923_398923;
   reg _398924_398924 ; 
   reg __398924_398924;
   reg _398925_398925 ; 
   reg __398925_398925;
   reg _398926_398926 ; 
   reg __398926_398926;
   reg _398927_398927 ; 
   reg __398927_398927;
   reg _398928_398928 ; 
   reg __398928_398928;
   reg _398929_398929 ; 
   reg __398929_398929;
   reg _398930_398930 ; 
   reg __398930_398930;
   reg _398931_398931 ; 
   reg __398931_398931;
   reg _398932_398932 ; 
   reg __398932_398932;
   reg _398933_398933 ; 
   reg __398933_398933;
   reg _398934_398934 ; 
   reg __398934_398934;
   reg _398935_398935 ; 
   reg __398935_398935;
   reg _398936_398936 ; 
   reg __398936_398936;
   reg _398937_398937 ; 
   reg __398937_398937;
   reg _398938_398938 ; 
   reg __398938_398938;
   reg _398939_398939 ; 
   reg __398939_398939;
   reg _398940_398940 ; 
   reg __398940_398940;
   reg _398941_398941 ; 
   reg __398941_398941;
   reg _398942_398942 ; 
   reg __398942_398942;
   reg _398943_398943 ; 
   reg __398943_398943;
   reg _398944_398944 ; 
   reg __398944_398944;
   reg _398945_398945 ; 
   reg __398945_398945;
   reg _398946_398946 ; 
   reg __398946_398946;
   reg _398947_398947 ; 
   reg __398947_398947;
   reg _398948_398948 ; 
   reg __398948_398948;
   reg _398949_398949 ; 
   reg __398949_398949;
   reg _398950_398950 ; 
   reg __398950_398950;
   reg _398951_398951 ; 
   reg __398951_398951;
   reg _398952_398952 ; 
   reg __398952_398952;
   reg _398953_398953 ; 
   reg __398953_398953;
   reg _398954_398954 ; 
   reg __398954_398954;
   reg _398955_398955 ; 
   reg __398955_398955;
   reg _398956_398956 ; 
   reg __398956_398956;
   reg _398957_398957 ; 
   reg __398957_398957;
   reg _398958_398958 ; 
   reg __398958_398958;
   reg _398959_398959 ; 
   reg __398959_398959;
   reg _398960_398960 ; 
   reg __398960_398960;
   reg _398961_398961 ; 
   reg __398961_398961;
   reg _398962_398962 ; 
   reg __398962_398962;
   reg _398963_398963 ; 
   reg __398963_398963;
   reg _398964_398964 ; 
   reg __398964_398964;
   reg _398965_398965 ; 
   reg __398965_398965;
   reg _398966_398966 ; 
   reg __398966_398966;
   reg _398967_398967 ; 
   reg __398967_398967;
   reg _398968_398968 ; 
   reg __398968_398968;
   reg _398969_398969 ; 
   reg __398969_398969;
   reg _398970_398970 ; 
   reg __398970_398970;
   reg _398971_398971 ; 
   reg __398971_398971;
   reg _398972_398972 ; 
   reg __398972_398972;
   reg _398973_398973 ; 
   reg __398973_398973;
   reg _398974_398974 ; 
   reg __398974_398974;
   reg _398975_398975 ; 
   reg __398975_398975;
   reg _398976_398976 ; 
   reg __398976_398976;
   reg _398977_398977 ; 
   reg __398977_398977;
   reg _398978_398978 ; 
   reg __398978_398978;
   reg _398979_398979 ; 
   reg __398979_398979;
   reg _398980_398980 ; 
   reg __398980_398980;
   reg _398981_398981 ; 
   reg __398981_398981;
   reg _398982_398982 ; 
   reg __398982_398982;
   reg _398983_398983 ; 
   reg __398983_398983;
   reg _398984_398984 ; 
   reg __398984_398984;
   reg _398985_398985 ; 
   reg __398985_398985;
   reg _398986_398986 ; 
   reg __398986_398986;
   reg _398987_398987 ; 
   reg __398987_398987;
   reg _398988_398988 ; 
   reg __398988_398988;
   reg _398989_398989 ; 
   reg __398989_398989;
   reg _398990_398990 ; 
   reg __398990_398990;
   reg _398991_398991 ; 
   reg __398991_398991;
   reg _398992_398992 ; 
   reg __398992_398992;
   reg _398993_398993 ; 
   reg __398993_398993;
   reg _398994_398994 ; 
   reg __398994_398994;
   reg _398995_398995 ; 
   reg __398995_398995;
   reg _398996_398996 ; 
   reg __398996_398996;
   reg _398997_398997 ; 
   reg __398997_398997;
   reg _398998_398998 ; 
   reg __398998_398998;
   reg _398999_398999 ; 
   reg __398999_398999;
   reg _399000_399000 ; 
   reg __399000_399000;
   reg _399001_399001 ; 
   reg __399001_399001;
   reg _399002_399002 ; 
   reg __399002_399002;
   reg _399003_399003 ; 
   reg __399003_399003;
   reg _399004_399004 ; 
   reg __399004_399004;
   reg _399005_399005 ; 
   reg __399005_399005;
   reg _399006_399006 ; 
   reg __399006_399006;
   reg _399007_399007 ; 
   reg __399007_399007;
   reg _399008_399008 ; 
   reg __399008_399008;
   reg _399009_399009 ; 
   reg __399009_399009;
   reg _399010_399010 ; 
   reg __399010_399010;
   reg _399011_399011 ; 
   reg __399011_399011;
   reg _399012_399012 ; 
   reg __399012_399012;
   reg _399013_399013 ; 
   reg __399013_399013;
   reg _399014_399014 ; 
   reg __399014_399014;
   reg _399015_399015 ; 
   reg __399015_399015;
   reg _399016_399016 ; 
   reg __399016_399016;
   reg _399017_399017 ; 
   reg __399017_399017;
   reg _399018_399018 ; 
   reg __399018_399018;
   reg _399019_399019 ; 
   reg __399019_399019;
   reg _399020_399020 ; 
   reg __399020_399020;
   reg _399021_399021 ; 
   reg __399021_399021;
   reg _399022_399022 ; 
   reg __399022_399022;
   reg _399023_399023 ; 
   reg __399023_399023;
   reg _399024_399024 ; 
   reg __399024_399024;
   reg _399025_399025 ; 
   reg __399025_399025;
   reg _399026_399026 ; 
   reg __399026_399026;
   reg _399027_399027 ; 
   reg __399027_399027;
   reg _399028_399028 ; 
   reg __399028_399028;
   reg _399029_399029 ; 
   reg __399029_399029;
   reg _399030_399030 ; 
   reg __399030_399030;
   reg _399031_399031 ; 
   reg __399031_399031;
   reg _399032_399032 ; 
   reg __399032_399032;
   reg _399033_399033 ; 
   reg __399033_399033;
   reg _399034_399034 ; 
   reg __399034_399034;
   reg _399035_399035 ; 
   reg __399035_399035;
   reg _399036_399036 ; 
   reg __399036_399036;
   reg _399037_399037 ; 
   reg __399037_399037;
   reg _399038_399038 ; 
   reg __399038_399038;
   reg _399039_399039 ; 
   reg __399039_399039;
   reg _399040_399040 ; 
   reg __399040_399040;
   reg _399041_399041 ; 
   reg __399041_399041;
   reg _399042_399042 ; 
   reg __399042_399042;
   reg _399043_399043 ; 
   reg __399043_399043;
   reg _399044_399044 ; 
   reg __399044_399044;
   reg _399045_399045 ; 
   reg __399045_399045;
   reg _399046_399046 ; 
   reg __399046_399046;
   reg _399047_399047 ; 
   reg __399047_399047;
   reg _399048_399048 ; 
   reg __399048_399048;
   reg _399049_399049 ; 
   reg __399049_399049;
   reg _399050_399050 ; 
   reg __399050_399050;
   reg _399051_399051 ; 
   reg __399051_399051;
   reg _399052_399052 ; 
   reg __399052_399052;
   reg _399053_399053 ; 
   reg __399053_399053;
   reg _399054_399054 ; 
   reg __399054_399054;
   reg _399055_399055 ; 
   reg __399055_399055;
   reg _399056_399056 ; 
   reg __399056_399056;
   reg _399057_399057 ; 
   reg __399057_399057;
   reg _399058_399058 ; 
   reg __399058_399058;
   reg _399059_399059 ; 
   reg __399059_399059;
   reg _399060_399060 ; 
   reg __399060_399060;
   reg _399061_399061 ; 
   reg __399061_399061;
   reg _399062_399062 ; 
   reg __399062_399062;
   reg _399063_399063 ; 
   reg __399063_399063;
   reg _399064_399064 ; 
   reg __399064_399064;
   reg _399065_399065 ; 
   reg __399065_399065;
   reg _399066_399066 ; 
   reg __399066_399066;
   reg _399067_399067 ; 
   reg __399067_399067;
   reg _399068_399068 ; 
   reg __399068_399068;
   reg _399069_399069 ; 
   reg __399069_399069;
   reg _399070_399070 ; 
   reg __399070_399070;
   reg _399071_399071 ; 
   reg __399071_399071;
   reg _399072_399072 ; 
   reg __399072_399072;
   reg _399073_399073 ; 
   reg __399073_399073;
   reg _399074_399074 ; 
   reg __399074_399074;
   reg _399075_399075 ; 
   reg __399075_399075;
   reg _399076_399076 ; 
   reg __399076_399076;
   reg _399077_399077 ; 
   reg __399077_399077;
   reg _399078_399078 ; 
   reg __399078_399078;
   reg _399079_399079 ; 
   reg __399079_399079;
   reg _399080_399080 ; 
   reg __399080_399080;
   reg _399081_399081 ; 
   reg __399081_399081;
   reg _399082_399082 ; 
   reg __399082_399082;
   reg _399083_399083 ; 
   reg __399083_399083;
   reg _399084_399084 ; 
   reg __399084_399084;
   reg _399085_399085 ; 
   reg __399085_399085;
   reg _399086_399086 ; 
   reg __399086_399086;
   reg _399087_399087 ; 
   reg __399087_399087;
   reg _399088_399088 ; 
   reg __399088_399088;
   reg _399089_399089 ; 
   reg __399089_399089;
   reg _399090_399090 ; 
   reg __399090_399090;
   reg _399091_399091 ; 
   reg __399091_399091;
   reg _399092_399092 ; 
   reg __399092_399092;
   reg _399093_399093 ; 
   reg __399093_399093;
   reg _399094_399094 ; 
   reg __399094_399094;
   reg _399095_399095 ; 
   reg __399095_399095;
   reg _399096_399096 ; 
   reg __399096_399096;
   reg _399097_399097 ; 
   reg __399097_399097;
   reg _399098_399098 ; 
   reg __399098_399098;
   reg _399099_399099 ; 
   reg __399099_399099;
   reg _399100_399100 ; 
   reg __399100_399100;
   reg _399101_399101 ; 
   reg __399101_399101;
   reg _399102_399102 ; 
   reg __399102_399102;
   reg _399103_399103 ; 
   reg __399103_399103;
   reg _399104_399104 ; 
   reg __399104_399104;
   reg _399105_399105 ; 
   reg __399105_399105;
   reg _399106_399106 ; 
   reg __399106_399106;
   reg _399107_399107 ; 
   reg __399107_399107;
   reg _399108_399108 ; 
   reg __399108_399108;
   reg _399109_399109 ; 
   reg __399109_399109;
   reg _399110_399110 ; 
   reg __399110_399110;
   reg _399111_399111 ; 
   reg __399111_399111;
   reg _399112_399112 ; 
   reg __399112_399112;
   reg _399113_399113 ; 
   reg __399113_399113;
   reg _399114_399114 ; 
   reg __399114_399114;
   reg _399115_399115 ; 
   reg __399115_399115;
   reg _399116_399116 ; 
   reg __399116_399116;
   reg _399117_399117 ; 
   reg __399117_399117;
   reg _399118_399118 ; 
   reg __399118_399118;
   reg _399119_399119 ; 
   reg __399119_399119;
   reg _399120_399120 ; 
   reg __399120_399120;
   reg _399121_399121 ; 
   reg __399121_399121;
   reg _399122_399122 ; 
   reg __399122_399122;
   reg _399123_399123 ; 
   reg __399123_399123;
   reg _399124_399124 ; 
   reg __399124_399124;
   reg _399125_399125 ; 
   reg __399125_399125;
   reg _399126_399126 ; 
   reg __399126_399126;
   reg _399127_399127 ; 
   reg __399127_399127;
   reg _399128_399128 ; 
   reg __399128_399128;
   reg _399129_399129 ; 
   reg __399129_399129;
   reg _399130_399130 ; 
   reg __399130_399130;
   reg _399131_399131 ; 
   reg __399131_399131;
   reg _399132_399132 ; 
   reg __399132_399132;
   reg _399133_399133 ; 
   reg __399133_399133;
   reg _399134_399134 ; 
   reg __399134_399134;
   reg _399135_399135 ; 
   reg __399135_399135;
   reg _399136_399136 ; 
   reg __399136_399136;
   reg _399137_399137 ; 
   reg __399137_399137;
   reg _399138_399138 ; 
   reg __399138_399138;
   reg _399139_399139 ; 
   reg __399139_399139;
   reg _399140_399140 ; 
   reg __399140_399140;
   reg _399141_399141 ; 
   reg __399141_399141;
   reg _399142_399142 ; 
   reg __399142_399142;
   reg _399143_399143 ; 
   reg __399143_399143;
   reg _399144_399144 ; 
   reg __399144_399144;
   reg _399145_399145 ; 
   reg __399145_399145;
   reg _399146_399146 ; 
   reg __399146_399146;
   reg _399147_399147 ; 
   reg __399147_399147;
   reg _399148_399148 ; 
   reg __399148_399148;
   reg _399149_399149 ; 
   reg __399149_399149;
   reg _399150_399150 ; 
   reg __399150_399150;
   reg _399151_399151 ; 
   reg __399151_399151;
   reg _399152_399152 ; 
   reg __399152_399152;
   reg _399153_399153 ; 
   reg __399153_399153;
   reg _399154_399154 ; 
   reg __399154_399154;
   reg _399155_399155 ; 
   reg __399155_399155;
   reg _399156_399156 ; 
   reg __399156_399156;
   reg _399157_399157 ; 
   reg __399157_399157;
   reg _399158_399158 ; 
   reg __399158_399158;
   reg _399159_399159 ; 
   reg __399159_399159;
   reg _399160_399160 ; 
   reg __399160_399160;
   reg _399161_399161 ; 
   reg __399161_399161;
   reg _399162_399162 ; 
   reg __399162_399162;
   reg _399163_399163 ; 
   reg __399163_399163;
   reg _399164_399164 ; 
   reg __399164_399164;
   reg _399165_399165 ; 
   reg __399165_399165;
   reg _399166_399166 ; 
   reg __399166_399166;
   reg _399167_399167 ; 
   reg __399167_399167;
   reg _399168_399168 ; 
   reg __399168_399168;
   reg _399169_399169 ; 
   reg __399169_399169;
   reg _399170_399170 ; 
   reg __399170_399170;
   reg _399171_399171 ; 
   reg __399171_399171;
   reg _399172_399172 ; 
   reg __399172_399172;
   reg _399173_399173 ; 
   reg __399173_399173;
   reg _399174_399174 ; 
   reg __399174_399174;
   reg _399175_399175 ; 
   reg __399175_399175;
   reg _399176_399176 ; 
   reg __399176_399176;
   reg _399177_399177 ; 
   reg __399177_399177;
   reg _399178_399178 ; 
   reg __399178_399178;
   reg _399179_399179 ; 
   reg __399179_399179;
   reg _399180_399180 ; 
   reg __399180_399180;
   reg _399181_399181 ; 
   reg __399181_399181;
   reg _399182_399182 ; 
   reg __399182_399182;
   reg _399183_399183 ; 
   reg __399183_399183;
   reg _399184_399184 ; 
   reg __399184_399184;
   reg _399185_399185 ; 
   reg __399185_399185;
   reg _399186_399186 ; 
   reg __399186_399186;
   reg _399187_399187 ; 
   reg __399187_399187;
   reg _399188_399188 ; 
   reg __399188_399188;
   reg _399189_399189 ; 
   reg __399189_399189;
   reg _399190_399190 ; 
   reg __399190_399190;
   reg _399191_399191 ; 
   reg __399191_399191;
   reg _399192_399192 ; 
   reg __399192_399192;
   reg _399193_399193 ; 
   reg __399193_399193;
   reg _399194_399194 ; 
   reg __399194_399194;
   reg _399195_399195 ; 
   reg __399195_399195;
   reg _399196_399196 ; 
   reg __399196_399196;
   reg _399197_399197 ; 
   reg __399197_399197;
   reg _399198_399198 ; 
   reg __399198_399198;
   reg _399199_399199 ; 
   reg __399199_399199;
   reg _399200_399200 ; 
   reg __399200_399200;
   reg _399201_399201 ; 
   reg __399201_399201;
   reg _399202_399202 ; 
   reg __399202_399202;
   reg _399203_399203 ; 
   reg __399203_399203;
   reg _399204_399204 ; 
   reg __399204_399204;
   reg _399205_399205 ; 
   reg __399205_399205;
   reg _399206_399206 ; 
   reg __399206_399206;
   reg _399207_399207 ; 
   reg __399207_399207;
   reg _399208_399208 ; 
   reg __399208_399208;
   reg _399209_399209 ; 
   reg __399209_399209;
   reg _399210_399210 ; 
   reg __399210_399210;
   reg _399211_399211 ; 
   reg __399211_399211;
   reg _399212_399212 ; 
   reg __399212_399212;
   reg _399213_399213 ; 
   reg __399213_399213;
   reg _399214_399214 ; 
   reg __399214_399214;
   reg _399215_399215 ; 
   reg __399215_399215;
   reg _399216_399216 ; 
   reg __399216_399216;
   reg _399217_399217 ; 
   reg __399217_399217;
   reg _399218_399218 ; 
   reg __399218_399218;
   reg _399219_399219 ; 
   reg __399219_399219;
   reg _399220_399220 ; 
   reg __399220_399220;
   reg _399221_399221 ; 
   reg __399221_399221;
   reg _399222_399222 ; 
   reg __399222_399222;
   reg _399223_399223 ; 
   reg __399223_399223;
   reg _399224_399224 ; 
   reg __399224_399224;
   reg _399225_399225 ; 
   reg __399225_399225;
   reg _399226_399226 ; 
   reg __399226_399226;
   reg _399227_399227 ; 
   reg __399227_399227;
   reg _399228_399228 ; 
   reg __399228_399228;
   reg _399229_399229 ; 
   reg __399229_399229;
   reg _399230_399230 ; 
   reg __399230_399230;
   reg _399231_399231 ; 
   reg __399231_399231;
   reg _399232_399232 ; 
   reg __399232_399232;
   reg _399233_399233 ; 
   reg __399233_399233;
   reg _399234_399234 ; 
   reg __399234_399234;
   reg _399235_399235 ; 
   reg __399235_399235;
   reg _399236_399236 ; 
   reg __399236_399236;
   reg _399237_399237 ; 
   reg __399237_399237;
   reg _399238_399238 ; 
   reg __399238_399238;
   reg _399239_399239 ; 
   reg __399239_399239;
   reg _399240_399240 ; 
   reg __399240_399240;
   reg _399241_399241 ; 
   reg __399241_399241;
   reg _399242_399242 ; 
   reg __399242_399242;
   reg _399243_399243 ; 
   reg __399243_399243;
   reg _399244_399244 ; 
   reg __399244_399244;
   reg _399245_399245 ; 
   reg __399245_399245;
   reg _399246_399246 ; 
   reg __399246_399246;
   reg _399247_399247 ; 
   reg __399247_399247;
   reg _399248_399248 ; 
   reg __399248_399248;
   reg _399249_399249 ; 
   reg __399249_399249;
   reg _399250_399250 ; 
   reg __399250_399250;
   reg _399251_399251 ; 
   reg __399251_399251;
   reg _399252_399252 ; 
   reg __399252_399252;
   reg _399253_399253 ; 
   reg __399253_399253;
   reg _399254_399254 ; 
   reg __399254_399254;
   reg _399255_399255 ; 
   reg __399255_399255;
   reg _399256_399256 ; 
   reg __399256_399256;
   reg _399257_399257 ; 
   reg __399257_399257;
   reg _399258_399258 ; 
   reg __399258_399258;
   reg _399259_399259 ; 
   reg __399259_399259;
   reg _399260_399260 ; 
   reg __399260_399260;
   reg _399261_399261 ; 
   reg __399261_399261;
   reg _399262_399262 ; 
   reg __399262_399262;
   reg _399263_399263 ; 
   reg __399263_399263;
   reg _399264_399264 ; 
   reg __399264_399264;
   reg _399265_399265 ; 
   reg __399265_399265;
   reg _399266_399266 ; 
   reg __399266_399266;
   reg _399267_399267 ; 
   reg __399267_399267;
   reg _399268_399268 ; 
   reg __399268_399268;
   reg _399269_399269 ; 
   reg __399269_399269;
   reg _399270_399270 ; 
   reg __399270_399270;
   reg _399271_399271 ; 
   reg __399271_399271;
   reg _399272_399272 ; 
   reg __399272_399272;
   reg _399273_399273 ; 
   reg __399273_399273;
   reg _399274_399274 ; 
   reg __399274_399274;
   reg _399275_399275 ; 
   reg __399275_399275;
   reg _399276_399276 ; 
   reg __399276_399276;
   reg _399277_399277 ; 
   reg __399277_399277;
   reg _399278_399278 ; 
   reg __399278_399278;
   reg _399279_399279 ; 
   reg __399279_399279;
   reg _399280_399280 ; 
   reg __399280_399280;
   reg _399281_399281 ; 
   reg __399281_399281;
   reg _399282_399282 ; 
   reg __399282_399282;
   reg _399283_399283 ; 
   reg __399283_399283;
   reg _399284_399284 ; 
   reg __399284_399284;
   reg _399285_399285 ; 
   reg __399285_399285;
   reg _399286_399286 ; 
   reg __399286_399286;
   reg _399287_399287 ; 
   reg __399287_399287;
   reg _399288_399288 ; 
   reg __399288_399288;
   reg _399289_399289 ; 
   reg __399289_399289;
   reg _399290_399290 ; 
   reg __399290_399290;
   reg _399291_399291 ; 
   reg __399291_399291;
   reg _399292_399292 ; 
   reg __399292_399292;
   reg _399293_399293 ; 
   reg __399293_399293;
   reg _399294_399294 ; 
   reg __399294_399294;
   reg _399295_399295 ; 
   reg __399295_399295;
   reg _399296_399296 ; 
   reg __399296_399296;
   reg _399297_399297 ; 
   reg __399297_399297;
   reg _399298_399298 ; 
   reg __399298_399298;
   reg _399299_399299 ; 
   reg __399299_399299;
   reg _399300_399300 ; 
   reg __399300_399300;
   reg _399301_399301 ; 
   reg __399301_399301;
   reg _399302_399302 ; 
   reg __399302_399302;
   reg _399303_399303 ; 
   reg __399303_399303;
   reg _399304_399304 ; 
   reg __399304_399304;
   reg _399305_399305 ; 
   reg __399305_399305;
   reg _399306_399306 ; 
   reg __399306_399306;
   reg _399307_399307 ; 
   reg __399307_399307;
   reg _399308_399308 ; 
   reg __399308_399308;
   reg _399309_399309 ; 
   reg __399309_399309;
   reg _399310_399310 ; 
   reg __399310_399310;
   reg _399311_399311 ; 
   reg __399311_399311;
   reg _399312_399312 ; 
   reg __399312_399312;
   reg _399313_399313 ; 
   reg __399313_399313;
   reg _399314_399314 ; 
   reg __399314_399314;
   reg _399315_399315 ; 
   reg __399315_399315;
   reg _399316_399316 ; 
   reg __399316_399316;
   reg _399317_399317 ; 
   reg __399317_399317;
   reg _399318_399318 ; 
   reg __399318_399318;
   reg _399319_399319 ; 
   reg __399319_399319;
   reg _399320_399320 ; 
   reg __399320_399320;
   reg _399321_399321 ; 
   reg __399321_399321;
   reg _399322_399322 ; 
   reg __399322_399322;
   reg _399323_399323 ; 
   reg __399323_399323;
   reg _399324_399324 ; 
   reg __399324_399324;
   reg _399325_399325 ; 
   reg __399325_399325;
   reg _399326_399326 ; 
   reg __399326_399326;
   reg _399327_399327 ; 
   reg __399327_399327;
   reg _399328_399328 ; 
   reg __399328_399328;
   reg _399329_399329 ; 
   reg __399329_399329;
   reg _399330_399330 ; 
   reg __399330_399330;
   reg _399331_399331 ; 
   reg __399331_399331;
   reg _399332_399332 ; 
   reg __399332_399332;
   reg _399333_399333 ; 
   reg __399333_399333;
   reg _399334_399334 ; 
   reg __399334_399334;
   reg _399335_399335 ; 
   reg __399335_399335;
   reg _399336_399336 ; 
   reg __399336_399336;
   reg _399337_399337 ; 
   reg __399337_399337;
   reg _399338_399338 ; 
   reg __399338_399338;
   reg _399339_399339 ; 
   reg __399339_399339;
   reg _399340_399340 ; 
   reg __399340_399340;
   reg _399341_399341 ; 
   reg __399341_399341;
   reg _399342_399342 ; 
   reg __399342_399342;
   reg _399343_399343 ; 
   reg __399343_399343;
   reg _399344_399344 ; 
   reg __399344_399344;
   reg _399345_399345 ; 
   reg __399345_399345;
   reg _399346_399346 ; 
   reg __399346_399346;
   reg _399347_399347 ; 
   reg __399347_399347;
   reg _399348_399348 ; 
   reg __399348_399348;
   reg _399349_399349 ; 
   reg __399349_399349;
   reg _399350_399350 ; 
   reg __399350_399350;
   reg _399351_399351 ; 
   reg __399351_399351;
   reg _399352_399352 ; 
   reg __399352_399352;
   reg _399353_399353 ; 
   reg __399353_399353;
   reg _399354_399354 ; 
   reg __399354_399354;
   reg _399355_399355 ; 
   reg __399355_399355;
   reg _399356_399356 ; 
   reg __399356_399356;
   reg _399357_399357 ; 
   reg __399357_399357;
   reg _399358_399358 ; 
   reg __399358_399358;
   reg _399359_399359 ; 
   reg __399359_399359;
   reg _399360_399360 ; 
   reg __399360_399360;
   reg _399361_399361 ; 
   reg __399361_399361;
   reg _399362_399362 ; 
   reg __399362_399362;
   reg _399363_399363 ; 
   reg __399363_399363;
   reg _399364_399364 ; 
   reg __399364_399364;
   reg _399365_399365 ; 
   reg __399365_399365;
   reg _399366_399366 ; 
   reg __399366_399366;
   reg _399367_399367 ; 
   reg __399367_399367;
   reg _399368_399368 ; 
   reg __399368_399368;
   reg _399369_399369 ; 
   reg __399369_399369;
   reg _399370_399370 ; 
   reg __399370_399370;
   reg _399371_399371 ; 
   reg __399371_399371;
   reg _399372_399372 ; 
   reg __399372_399372;
   reg _399373_399373 ; 
   reg __399373_399373;
   reg _399374_399374 ; 
   reg __399374_399374;
   reg _399375_399375 ; 
   reg __399375_399375;
   reg _399376_399376 ; 
   reg __399376_399376;
   reg _399377_399377 ; 
   reg __399377_399377;
   reg _399378_399378 ; 
   reg __399378_399378;
   reg _399379_399379 ; 
   reg __399379_399379;
   reg _399380_399380 ; 
   reg __399380_399380;
   reg _399381_399381 ; 
   reg __399381_399381;
   reg _399382_399382 ; 
   reg __399382_399382;
   reg _399383_399383 ; 
   reg __399383_399383;
   reg _399384_399384 ; 
   reg __399384_399384;
   reg _399385_399385 ; 
   reg __399385_399385;
   reg _399386_399386 ; 
   reg __399386_399386;
   reg _399387_399387 ; 
   reg __399387_399387;
   reg _399388_399388 ; 
   reg __399388_399388;
   reg _399389_399389 ; 
   reg __399389_399389;
   reg _399390_399390 ; 
   reg __399390_399390;
   reg _399391_399391 ; 
   reg __399391_399391;
   reg _399392_399392 ; 
   reg __399392_399392;
   reg _399393_399393 ; 
   reg __399393_399393;
   reg _399394_399394 ; 
   reg __399394_399394;
   reg _399395_399395 ; 
   reg __399395_399395;
   reg _399396_399396 ; 
   reg __399396_399396;
   reg _399397_399397 ; 
   reg __399397_399397;
   reg _399398_399398 ; 
   reg __399398_399398;
   reg _399399_399399 ; 
   reg __399399_399399;
   reg _399400_399400 ; 
   reg __399400_399400;
   reg _399401_399401 ; 
   reg __399401_399401;
   reg _399402_399402 ; 
   reg __399402_399402;
   reg _399403_399403 ; 
   reg __399403_399403;
   reg _399404_399404 ; 
   reg __399404_399404;
   reg _399405_399405 ; 
   reg __399405_399405;
   reg _399406_399406 ; 
   reg __399406_399406;
   reg _399407_399407 ; 
   reg __399407_399407;
   reg _399408_399408 ; 
   reg __399408_399408;
   reg _399409_399409 ; 
   reg __399409_399409;
   reg _399410_399410 ; 
   reg __399410_399410;
   reg _399411_399411 ; 
   reg __399411_399411;
   reg _399412_399412 ; 
   reg __399412_399412;
   reg _399413_399413 ; 
   reg __399413_399413;
   reg _399414_399414 ; 
   reg __399414_399414;
   reg _399415_399415 ; 
   reg __399415_399415;
   reg _399416_399416 ; 
   reg __399416_399416;
   reg _399417_399417 ; 
   reg __399417_399417;
   reg _399418_399418 ; 
   reg __399418_399418;
   reg _399419_399419 ; 
   reg __399419_399419;
   reg _399420_399420 ; 
   reg __399420_399420;
   reg _399421_399421 ; 
   reg __399421_399421;
   reg _399422_399422 ; 
   reg __399422_399422;
   reg _399423_399423 ; 
   reg __399423_399423;
   reg _399424_399424 ; 
   reg __399424_399424;
   reg _399425_399425 ; 
   reg __399425_399425;
   reg _399426_399426 ; 
   reg __399426_399426;
   reg _399427_399427 ; 
   reg __399427_399427;
   reg _399428_399428 ; 
   reg __399428_399428;
   reg _399429_399429 ; 
   reg __399429_399429;
   reg _399430_399430 ; 
   reg __399430_399430;
   reg _399431_399431 ; 
   reg __399431_399431;
   reg _399432_399432 ; 
   reg __399432_399432;
   reg _399433_399433 ; 
   reg __399433_399433;
   reg _399434_399434 ; 
   reg __399434_399434;
   reg _399435_399435 ; 
   reg __399435_399435;
   reg _399436_399436 ; 
   reg __399436_399436;
   reg _399437_399437 ; 
   reg __399437_399437;
   reg _399438_399438 ; 
   reg __399438_399438;
   reg _399439_399439 ; 
   reg __399439_399439;
   reg _399440_399440 ; 
   reg __399440_399440;
   reg _399441_399441 ; 
   reg __399441_399441;
   reg _399442_399442 ; 
   reg __399442_399442;
   reg _399443_399443 ; 
   reg __399443_399443;
   reg _399444_399444 ; 
   reg __399444_399444;
   reg _399445_399445 ; 
   reg __399445_399445;
   reg _399446_399446 ; 
   reg __399446_399446;
   reg _399447_399447 ; 
   reg __399447_399447;
   reg _399448_399448 ; 
   reg __399448_399448;
   reg _399449_399449 ; 
   reg __399449_399449;
   reg _399450_399450 ; 
   reg __399450_399450;
   reg _399451_399451 ; 
   reg __399451_399451;
   reg _399452_399452 ; 
   reg __399452_399452;
   reg _399453_399453 ; 
   reg __399453_399453;
   reg _399454_399454 ; 
   reg __399454_399454;
   reg _399455_399455 ; 
   reg __399455_399455;
   reg _399456_399456 ; 
   reg __399456_399456;
   reg _399457_399457 ; 
   reg __399457_399457;
   reg _399458_399458 ; 
   reg __399458_399458;
   reg _399459_399459 ; 
   reg __399459_399459;
   reg _399460_399460 ; 
   reg __399460_399460;
   reg _399461_399461 ; 
   reg __399461_399461;
   reg _399462_399462 ; 
   reg __399462_399462;
   reg _399463_399463 ; 
   reg __399463_399463;
   reg _399464_399464 ; 
   reg __399464_399464;
   reg _399465_399465 ; 
   reg __399465_399465;
   reg _399466_399466 ; 
   reg __399466_399466;
   reg _399467_399467 ; 
   reg __399467_399467;
   reg _399468_399468 ; 
   reg __399468_399468;
   reg _399469_399469 ; 
   reg __399469_399469;
   reg _399470_399470 ; 
   reg __399470_399470;
   reg _399471_399471 ; 
   reg __399471_399471;
   reg _399472_399472 ; 
   reg __399472_399472;
   reg _399473_399473 ; 
   reg __399473_399473;
   reg _399474_399474 ; 
   reg __399474_399474;
   reg _399475_399475 ; 
   reg __399475_399475;
   reg _399476_399476 ; 
   reg __399476_399476;
   reg _399477_399477 ; 
   reg __399477_399477;
   reg _399478_399478 ; 
   reg __399478_399478;
   reg _399479_399479 ; 
   reg __399479_399479;
   reg _399480_399480 ; 
   reg __399480_399480;
   reg _399481_399481 ; 
   reg __399481_399481;
   reg _399482_399482 ; 
   reg __399482_399482;
   reg _399483_399483 ; 
   reg __399483_399483;
   reg _399484_399484 ; 
   reg __399484_399484;
   reg _399485_399485 ; 
   reg __399485_399485;
   reg _399486_399486 ; 
   reg __399486_399486;
   reg _399487_399487 ; 
   reg __399487_399487;
   reg _399488_399488 ; 
   reg __399488_399488;
   reg _399489_399489 ; 
   reg __399489_399489;
   reg _399490_399490 ; 
   reg __399490_399490;
   reg _399491_399491 ; 
   reg __399491_399491;
   reg _399492_399492 ; 
   reg __399492_399492;
   reg _399493_399493 ; 
   reg __399493_399493;
   reg _399494_399494 ; 
   reg __399494_399494;
   reg _399495_399495 ; 
   reg __399495_399495;
   reg _399496_399496 ; 
   reg __399496_399496;
   reg _399497_399497 ; 
   reg __399497_399497;
   reg _399498_399498 ; 
   reg __399498_399498;
   reg _399499_399499 ; 
   reg __399499_399499;
   reg _399500_399500 ; 
   reg __399500_399500;
   reg _399501_399501 ; 
   reg __399501_399501;
   reg _399502_399502 ; 
   reg __399502_399502;
   reg _399503_399503 ; 
   reg __399503_399503;
   reg _399504_399504 ; 
   reg __399504_399504;
   reg _399505_399505 ; 
   reg __399505_399505;
   reg _399506_399506 ; 
   reg __399506_399506;
   reg _399507_399507 ; 
   reg __399507_399507;
   reg _399508_399508 ; 
   reg __399508_399508;
   reg _399509_399509 ; 
   reg __399509_399509;
   reg _399510_399510 ; 
   reg __399510_399510;
   reg _399511_399511 ; 
   reg __399511_399511;
   reg _399512_399512 ; 
   reg __399512_399512;
   reg _399513_399513 ; 
   reg __399513_399513;
   reg _399514_399514 ; 
   reg __399514_399514;
   reg _399515_399515 ; 
   reg __399515_399515;
   reg _399516_399516 ; 
   reg __399516_399516;
   reg _399517_399517 ; 
   reg __399517_399517;
   reg _399518_399518 ; 
   reg __399518_399518;
   reg _399519_399519 ; 
   reg __399519_399519;
   reg _399520_399520 ; 
   reg __399520_399520;
   reg _399521_399521 ; 
   reg __399521_399521;
   reg _399522_399522 ; 
   reg __399522_399522;
   reg _399523_399523 ; 
   reg __399523_399523;
   reg _399524_399524 ; 
   reg __399524_399524;
   reg _399525_399525 ; 
   reg __399525_399525;
   reg _399526_399526 ; 
   reg __399526_399526;
   reg _399527_399527 ; 
   reg __399527_399527;
   reg _399528_399528 ; 
   reg __399528_399528;
   reg _399529_399529 ; 
   reg __399529_399529;
   reg _399530_399530 ; 
   reg __399530_399530;
   reg _399531_399531 ; 
   reg __399531_399531;
   reg _399532_399532 ; 
   reg __399532_399532;
   reg _399533_399533 ; 
   reg __399533_399533;
   reg _399534_399534 ; 
   reg __399534_399534;
   reg _399535_399535 ; 
   reg __399535_399535;
   reg _399536_399536 ; 
   reg __399536_399536;
   reg _399537_399537 ; 
   reg __399537_399537;
   reg _399538_399538 ; 
   reg __399538_399538;
   reg _399539_399539 ; 
   reg __399539_399539;
   reg _399540_399540 ; 
   reg __399540_399540;
   reg _399541_399541 ; 
   reg __399541_399541;
   reg _399542_399542 ; 
   reg __399542_399542;
   reg _399543_399543 ; 
   reg __399543_399543;
   reg _399544_399544 ; 
   reg __399544_399544;
   reg _399545_399545 ; 
   reg __399545_399545;
   reg _399546_399546 ; 
   reg __399546_399546;
   reg _399547_399547 ; 
   reg __399547_399547;
   reg _399548_399548 ; 
   reg __399548_399548;
   reg _399549_399549 ; 
   reg __399549_399549;
   reg _399550_399550 ; 
   reg __399550_399550;
   reg _399551_399551 ; 
   reg __399551_399551;
   reg _399552_399552 ; 
   reg __399552_399552;
   reg _399553_399553 ; 
   reg __399553_399553;
   reg _399554_399554 ; 
   reg __399554_399554;
   reg _399555_399555 ; 
   reg __399555_399555;
   reg _399556_399556 ; 
   reg __399556_399556;
   reg _399557_399557 ; 
   reg __399557_399557;
   reg _399558_399558 ; 
   reg __399558_399558;
   reg _399559_399559 ; 
   reg __399559_399559;
   reg _399560_399560 ; 
   reg __399560_399560;
   reg _399561_399561 ; 
   reg __399561_399561;
   reg _399562_399562 ; 
   reg __399562_399562;
   reg _399563_399563 ; 
   reg __399563_399563;
   reg _399564_399564 ; 
   reg __399564_399564;
   reg _399565_399565 ; 
   reg __399565_399565;
   reg _399566_399566 ; 
   reg __399566_399566;
   reg _399567_399567 ; 
   reg __399567_399567;
   reg _399568_399568 ; 
   reg __399568_399568;
   reg _399569_399569 ; 
   reg __399569_399569;
   reg _399570_399570 ; 
   reg __399570_399570;
   reg _399571_399571 ; 
   reg __399571_399571;
   reg _399572_399572 ; 
   reg __399572_399572;
   reg _399573_399573 ; 
   reg __399573_399573;
   reg _399574_399574 ; 
   reg __399574_399574;
   reg _399575_399575 ; 
   reg __399575_399575;
   reg _399576_399576 ; 
   reg __399576_399576;
   reg _399577_399577 ; 
   reg __399577_399577;
   reg _399578_399578 ; 
   reg __399578_399578;
   reg _399579_399579 ; 
   reg __399579_399579;
   reg _399580_399580 ; 
   reg __399580_399580;
   reg _399581_399581 ; 
   reg __399581_399581;
   reg _399582_399582 ; 
   reg __399582_399582;
   reg _399583_399583 ; 
   reg __399583_399583;
   reg _399584_399584 ; 
   reg __399584_399584;
   reg _399585_399585 ; 
   reg __399585_399585;
   reg _399586_399586 ; 
   reg __399586_399586;
   reg _399587_399587 ; 
   reg __399587_399587;
   reg _399588_399588 ; 
   reg __399588_399588;
   reg _399589_399589 ; 
   reg __399589_399589;
   reg _399590_399590 ; 
   reg __399590_399590;
   reg _399591_399591 ; 
   reg __399591_399591;
   reg _399592_399592 ; 
   reg __399592_399592;
   reg _399593_399593 ; 
   reg __399593_399593;
   reg _399594_399594 ; 
   reg __399594_399594;
   reg _399595_399595 ; 
   reg __399595_399595;
   reg _399596_399596 ; 
   reg __399596_399596;
   reg _399597_399597 ; 
   reg __399597_399597;
   reg _399598_399598 ; 
   reg __399598_399598;
   reg _399599_399599 ; 
   reg __399599_399599;
   reg _399600_399600 ; 
   reg __399600_399600;
   reg _399601_399601 ; 
   reg __399601_399601;
   reg _399602_399602 ; 
   reg __399602_399602;
   reg _399603_399603 ; 
   reg __399603_399603;
   reg _399604_399604 ; 
   reg __399604_399604;
   reg _399605_399605 ; 
   reg __399605_399605;
   reg _399606_399606 ; 
   reg __399606_399606;
   reg _399607_399607 ; 
   reg __399607_399607;
   reg _399608_399608 ; 
   reg __399608_399608;
   reg _399609_399609 ; 
   reg __399609_399609;
   reg _399610_399610 ; 
   reg __399610_399610;
   reg _399611_399611 ; 
   reg __399611_399611;
   reg _399612_399612 ; 
   reg __399612_399612;
   reg _399613_399613 ; 
   reg __399613_399613;
   reg _399614_399614 ; 
   reg __399614_399614;
   reg _399615_399615 ; 
   reg __399615_399615;
   reg _399616_399616 ; 
   reg __399616_399616;
   reg _399617_399617 ; 
   reg __399617_399617;
   reg _399618_399618 ; 
   reg __399618_399618;
   reg _399619_399619 ; 
   reg __399619_399619;
   reg _399620_399620 ; 
   reg __399620_399620;
   reg _399621_399621 ; 
   reg __399621_399621;
   reg _399622_399622 ; 
   reg __399622_399622;
   reg _399623_399623 ; 
   reg __399623_399623;
   reg _399624_399624 ; 
   reg __399624_399624;
   reg _399625_399625 ; 
   reg __399625_399625;
   reg _399626_399626 ; 
   reg __399626_399626;
   reg _399627_399627 ; 
   reg __399627_399627;
   reg _399628_399628 ; 
   reg __399628_399628;
   reg _399629_399629 ; 
   reg __399629_399629;
   reg _399630_399630 ; 
   reg __399630_399630;
   reg _399631_399631 ; 
   reg __399631_399631;
   reg _399632_399632 ; 
   reg __399632_399632;
   reg _399633_399633 ; 
   reg __399633_399633;
   reg _399634_399634 ; 
   reg __399634_399634;
   reg _399635_399635 ; 
   reg __399635_399635;
   reg _399636_399636 ; 
   reg __399636_399636;
   reg _399637_399637 ; 
   reg __399637_399637;
   reg _399638_399638 ; 
   reg __399638_399638;
   reg _399639_399639 ; 
   reg __399639_399639;
   reg _399640_399640 ; 
   reg __399640_399640;
   reg _399641_399641 ; 
   reg __399641_399641;
   reg _399642_399642 ; 
   reg __399642_399642;
   reg _399643_399643 ; 
   reg __399643_399643;
   reg _399644_399644 ; 
   reg __399644_399644;
   reg _399645_399645 ; 
   reg __399645_399645;
   reg _399646_399646 ; 
   reg __399646_399646;
   reg _399647_399647 ; 
   reg __399647_399647;
   reg _399648_399648 ; 
   reg __399648_399648;
   reg _399649_399649 ; 
   reg __399649_399649;
   reg _399650_399650 ; 
   reg __399650_399650;
   reg _399651_399651 ; 
   reg __399651_399651;
   reg _399652_399652 ; 
   reg __399652_399652;
   reg _399653_399653 ; 
   reg __399653_399653;
   reg _399654_399654 ; 
   reg __399654_399654;
   reg _399655_399655 ; 
   reg __399655_399655;
   reg _399656_399656 ; 
   reg __399656_399656;
   reg _399657_399657 ; 
   reg __399657_399657;
   reg _399658_399658 ; 
   reg __399658_399658;
   reg _399659_399659 ; 
   reg __399659_399659;
   reg _399660_399660 ; 
   reg __399660_399660;
   reg _399661_399661 ; 
   reg __399661_399661;
   reg _399662_399662 ; 
   reg __399662_399662;
   reg _399663_399663 ; 
   reg __399663_399663;
   reg _399664_399664 ; 
   reg __399664_399664;
   reg _399665_399665 ; 
   reg __399665_399665;
   reg _399666_399666 ; 
   reg __399666_399666;
   reg _399667_399667 ; 
   reg __399667_399667;
   reg _399668_399668 ; 
   reg __399668_399668;
   reg _399669_399669 ; 
   reg __399669_399669;
   reg _399670_399670 ; 
   reg __399670_399670;
   reg _399671_399671 ; 
   reg __399671_399671;
   reg _399672_399672 ; 
   reg __399672_399672;
   reg _399673_399673 ; 
   reg __399673_399673;
   reg _399674_399674 ; 
   reg __399674_399674;
   reg _399675_399675 ; 
   reg __399675_399675;
   reg _399676_399676 ; 
   reg __399676_399676;
   reg _399677_399677 ; 
   reg __399677_399677;
   reg _399678_399678 ; 
   reg __399678_399678;
   reg _399679_399679 ; 
   reg __399679_399679;
   reg _399680_399680 ; 
   reg __399680_399680;
   reg _399681_399681 ; 
   reg __399681_399681;
   reg _399682_399682 ; 
   reg __399682_399682;
   reg _399683_399683 ; 
   reg __399683_399683;
   reg _399684_399684 ; 
   reg __399684_399684;
   reg _399685_399685 ; 
   reg __399685_399685;
   reg _399686_399686 ; 
   reg __399686_399686;
   reg _399687_399687 ; 
   reg __399687_399687;
   reg _399688_399688 ; 
   reg __399688_399688;
   reg _399689_399689 ; 
   reg __399689_399689;
   reg _399690_399690 ; 
   reg __399690_399690;
   reg _399691_399691 ; 
   reg __399691_399691;
   reg _399692_399692 ; 
   reg __399692_399692;
   reg _399693_399693 ; 
   reg __399693_399693;
   reg _399694_399694 ; 
   reg __399694_399694;
   reg _399695_399695 ; 
   reg __399695_399695;
   reg _399696_399696 ; 
   reg __399696_399696;
   reg _399697_399697 ; 
   reg __399697_399697;
   reg _399698_399698 ; 
   reg __399698_399698;
   reg _399699_399699 ; 
   reg __399699_399699;
   reg _399700_399700 ; 
   reg __399700_399700;
   reg _399701_399701 ; 
   reg __399701_399701;
   reg _399702_399702 ; 
   reg __399702_399702;
   reg _399703_399703 ; 
   reg __399703_399703;
   reg _399704_399704 ; 
   reg __399704_399704;
   reg _399705_399705 ; 
   reg __399705_399705;
   reg _399706_399706 ; 
   reg __399706_399706;
   reg _399707_399707 ; 
   reg __399707_399707;
   reg _399708_399708 ; 
   reg __399708_399708;
   reg _399709_399709 ; 
   reg __399709_399709;
   reg _399710_399710 ; 
   reg __399710_399710;
   reg _399711_399711 ; 
   reg __399711_399711;
   reg _399712_399712 ; 
   reg __399712_399712;
   reg _399713_399713 ; 
   reg __399713_399713;
   reg _399714_399714 ; 
   reg __399714_399714;
   reg _399715_399715 ; 
   reg __399715_399715;
   reg _399716_399716 ; 
   reg __399716_399716;
   reg _399717_399717 ; 
   reg __399717_399717;
   reg _399718_399718 ; 
   reg __399718_399718;
   reg _399719_399719 ; 
   reg __399719_399719;
   reg _399720_399720 ; 
   reg __399720_399720;
   reg _399721_399721 ; 
   reg __399721_399721;
   reg _399722_399722 ; 
   reg __399722_399722;
   reg _399723_399723 ; 
   reg __399723_399723;
   reg _399724_399724 ; 
   reg __399724_399724;
   reg _399725_399725 ; 
   reg __399725_399725;
   reg _399726_399726 ; 
   reg __399726_399726;
   reg _399727_399727 ; 
   reg __399727_399727;
   reg _399728_399728 ; 
   reg __399728_399728;
   reg _399729_399729 ; 
   reg __399729_399729;
   reg _399730_399730 ; 
   reg __399730_399730;
   reg _399731_399731 ; 
   reg __399731_399731;
   reg _399732_399732 ; 
   reg __399732_399732;
   reg _399733_399733 ; 
   reg __399733_399733;
   reg _399734_399734 ; 
   reg __399734_399734;
   reg _399735_399735 ; 
   reg __399735_399735;
   reg _399736_399736 ; 
   reg __399736_399736;
   reg _399737_399737 ; 
   reg __399737_399737;
   reg _399738_399738 ; 
   reg __399738_399738;
   reg _399739_399739 ; 
   reg __399739_399739;
   reg _399740_399740 ; 
   reg __399740_399740;
   reg _399741_399741 ; 
   reg __399741_399741;
   reg _399742_399742 ; 
   reg __399742_399742;
   reg _399743_399743 ; 
   reg __399743_399743;
   reg _399744_399744 ; 
   reg __399744_399744;
   reg _399745_399745 ; 
   reg __399745_399745;
   reg _399746_399746 ; 
   reg __399746_399746;
   reg _399747_399747 ; 
   reg __399747_399747;
   reg _399748_399748 ; 
   reg __399748_399748;
   reg _399749_399749 ; 
   reg __399749_399749;
   reg _399750_399750 ; 
   reg __399750_399750;
   reg _399751_399751 ; 
   reg __399751_399751;
   reg _399752_399752 ; 
   reg __399752_399752;
   reg _399753_399753 ; 
   reg __399753_399753;
   reg _399754_399754 ; 
   reg __399754_399754;
   reg _399755_399755 ; 
   reg __399755_399755;
   reg _399756_399756 ; 
   reg __399756_399756;
   reg _399757_399757 ; 
   reg __399757_399757;
   reg _399758_399758 ; 
   reg __399758_399758;
   reg _399759_399759 ; 
   reg __399759_399759;
   reg _399760_399760 ; 
   reg __399760_399760;
   reg _399761_399761 ; 
   reg __399761_399761;
   reg _399762_399762 ; 
   reg __399762_399762;
   reg _399763_399763 ; 
   reg __399763_399763;
   reg _399764_399764 ; 
   reg __399764_399764;
   reg _399765_399765 ; 
   reg __399765_399765;
   reg _399766_399766 ; 
   reg __399766_399766;
   reg _399767_399767 ; 
   reg __399767_399767;
   reg _399768_399768 ; 
   reg __399768_399768;
   reg _399769_399769 ; 
   reg __399769_399769;
   reg _399770_399770 ; 
   reg __399770_399770;
   reg _399771_399771 ; 
   reg __399771_399771;
   reg _399772_399772 ; 
   reg __399772_399772;
   reg _399773_399773 ; 
   reg __399773_399773;
   reg _399774_399774 ; 
   reg __399774_399774;
   reg _399775_399775 ; 
   reg __399775_399775;
   reg _399776_399776 ; 
   reg __399776_399776;
   reg _399777_399777 ; 
   reg __399777_399777;
   reg _399778_399778 ; 
   reg __399778_399778;
   reg _399779_399779 ; 
   reg __399779_399779;
   reg _399780_399780 ; 
   reg __399780_399780;
   reg _399781_399781 ; 
   reg __399781_399781;
   reg _399782_399782 ; 
   reg __399782_399782;
   reg _399783_399783 ; 
   reg __399783_399783;
   reg _399784_399784 ; 
   reg __399784_399784;
   reg _399785_399785 ; 
   reg __399785_399785;
   reg _399786_399786 ; 
   reg __399786_399786;
   reg _399787_399787 ; 
   reg __399787_399787;
   reg _399788_399788 ; 
   reg __399788_399788;
   reg _399789_399789 ; 
   reg __399789_399789;
   reg _399790_399790 ; 
   reg __399790_399790;
   reg _399791_399791 ; 
   reg __399791_399791;
   reg _399792_399792 ; 
   reg __399792_399792;
   reg _399793_399793 ; 
   reg __399793_399793;
   reg _399794_399794 ; 
   reg __399794_399794;
   reg _399795_399795 ; 
   reg __399795_399795;
   reg _399796_399796 ; 
   reg __399796_399796;
   reg _399797_399797 ; 
   reg __399797_399797;
   reg _399798_399798 ; 
   reg __399798_399798;
   reg _399799_399799 ; 
   reg __399799_399799;
   reg _399800_399800 ; 
   reg __399800_399800;
   reg _399801_399801 ; 
   reg __399801_399801;
   reg _399802_399802 ; 
   reg __399802_399802;
   reg _399803_399803 ; 
   reg __399803_399803;
   reg _399804_399804 ; 
   reg __399804_399804;
   reg _399805_399805 ; 
   reg __399805_399805;
   reg _399806_399806 ; 
   reg __399806_399806;
   reg _399807_399807 ; 
   reg __399807_399807;
   reg _399808_399808 ; 
   reg __399808_399808;
   reg _399809_399809 ; 
   reg __399809_399809;
   reg _399810_399810 ; 
   reg __399810_399810;
   reg _399811_399811 ; 
   reg __399811_399811;
   reg _399812_399812 ; 
   reg __399812_399812;
   reg _399813_399813 ; 
   reg __399813_399813;
   reg _399814_399814 ; 
   reg __399814_399814;
   reg _399815_399815 ; 
   reg __399815_399815;
   reg _399816_399816 ; 
   reg __399816_399816;
   reg _399817_399817 ; 
   reg __399817_399817;
   reg _399818_399818 ; 
   reg __399818_399818;
   reg _399819_399819 ; 
   reg __399819_399819;
   reg _399820_399820 ; 
   reg __399820_399820;
   reg _399821_399821 ; 
   reg __399821_399821;
   reg _399822_399822 ; 
   reg __399822_399822;
   reg _399823_399823 ; 
   reg __399823_399823;
   reg _399824_399824 ; 
   reg __399824_399824;
   reg _399825_399825 ; 
   reg __399825_399825;
   reg _399826_399826 ; 
   reg __399826_399826;
   reg _399827_399827 ; 
   reg __399827_399827;
   reg _399828_399828 ; 
   reg __399828_399828;
   reg _399829_399829 ; 
   reg __399829_399829;
   reg _399830_399830 ; 
   reg __399830_399830;
   reg _399831_399831 ; 
   reg __399831_399831;
   reg _399832_399832 ; 
   reg __399832_399832;
   reg _399833_399833 ; 
   reg __399833_399833;
   reg _399834_399834 ; 
   reg __399834_399834;
   reg _399835_399835 ; 
   reg __399835_399835;
   reg _399836_399836 ; 
   reg __399836_399836;
   reg _399837_399837 ; 
   reg __399837_399837;
   reg _399838_399838 ; 
   reg __399838_399838;
   reg _399839_399839 ; 
   reg __399839_399839;
   reg _399840_399840 ; 
   reg __399840_399840;
   reg _399841_399841 ; 
   reg __399841_399841;
   reg _399842_399842 ; 
   reg __399842_399842;
   reg _399843_399843 ; 
   reg __399843_399843;
   reg _399844_399844 ; 
   reg __399844_399844;
   reg _399845_399845 ; 
   reg __399845_399845;
   reg _399846_399846 ; 
   reg __399846_399846;
   reg _399847_399847 ; 
   reg __399847_399847;
   reg _399848_399848 ; 
   reg __399848_399848;
   reg _399849_399849 ; 
   reg __399849_399849;
   reg _399850_399850 ; 
   reg __399850_399850;
   reg _399851_399851 ; 
   reg __399851_399851;
   reg _399852_399852 ; 
   reg __399852_399852;
   reg _399853_399853 ; 
   reg __399853_399853;
   reg _399854_399854 ; 
   reg __399854_399854;
   reg _399855_399855 ; 
   reg __399855_399855;
   reg _399856_399856 ; 
   reg __399856_399856;
   reg _399857_399857 ; 
   reg __399857_399857;
   reg _399858_399858 ; 
   reg __399858_399858;
   reg _399859_399859 ; 
   reg __399859_399859;
   reg _399860_399860 ; 
   reg __399860_399860;
   reg _399861_399861 ; 
   reg __399861_399861;
   reg _399862_399862 ; 
   reg __399862_399862;
   reg _399863_399863 ; 
   reg __399863_399863;
   reg _399864_399864 ; 
   reg __399864_399864;
   reg _399865_399865 ; 
   reg __399865_399865;
   reg _399866_399866 ; 
   reg __399866_399866;
   reg _399867_399867 ; 
   reg __399867_399867;
   reg _399868_399868 ; 
   reg __399868_399868;
   reg _399869_399869 ; 
   reg __399869_399869;
   reg _399870_399870 ; 
   reg __399870_399870;
   reg _399871_399871 ; 
   reg __399871_399871;
   reg _399872_399872 ; 
   reg __399872_399872;
   reg _399873_399873 ; 
   reg __399873_399873;
   reg _399874_399874 ; 
   reg __399874_399874;
   reg _399875_399875 ; 
   reg __399875_399875;
   reg _399876_399876 ; 
   reg __399876_399876;
   reg _399877_399877 ; 
   reg __399877_399877;
   reg _399878_399878 ; 
   reg __399878_399878;
   reg _399879_399879 ; 
   reg __399879_399879;
   reg _399880_399880 ; 
   reg __399880_399880;
   reg _399881_399881 ; 
   reg __399881_399881;
   reg _399882_399882 ; 
   reg __399882_399882;
   reg _399883_399883 ; 
   reg __399883_399883;
   reg _399884_399884 ; 
   reg __399884_399884;
   reg _399885_399885 ; 
   reg __399885_399885;
   reg _399886_399886 ; 
   reg __399886_399886;
   reg _399887_399887 ; 
   reg __399887_399887;
   reg _399888_399888 ; 
   reg __399888_399888;
   reg _399889_399889 ; 
   reg __399889_399889;
   reg _399890_399890 ; 
   reg __399890_399890;
   reg _399891_399891 ; 
   reg __399891_399891;
   reg _399892_399892 ; 
   reg __399892_399892;
   reg _399893_399893 ; 
   reg __399893_399893;
   reg _399894_399894 ; 
   reg __399894_399894;
   reg _399895_399895 ; 
   reg __399895_399895;
   reg _399896_399896 ; 
   reg __399896_399896;
   reg _399897_399897 ; 
   reg __399897_399897;
   reg _399898_399898 ; 
   reg __399898_399898;
   reg _399899_399899 ; 
   reg __399899_399899;
   reg _399900_399900 ; 
   reg __399900_399900;
   reg _399901_399901 ; 
   reg __399901_399901;
   reg _399902_399902 ; 
   reg __399902_399902;
   reg _399903_399903 ; 
   reg __399903_399903;
   reg _399904_399904 ; 
   reg __399904_399904;
   reg _399905_399905 ; 
   reg __399905_399905;
   reg _399906_399906 ; 
   reg __399906_399906;
   reg _399907_399907 ; 
   reg __399907_399907;
   reg _399908_399908 ; 
   reg __399908_399908;
   reg _399909_399909 ; 
   reg __399909_399909;
   reg _399910_399910 ; 
   reg __399910_399910;
   reg _399911_399911 ; 
   reg __399911_399911;
   reg _399912_399912 ; 
   reg __399912_399912;
   reg _399913_399913 ; 
   reg __399913_399913;
   reg _399914_399914 ; 
   reg __399914_399914;
   reg _399915_399915 ; 
   reg __399915_399915;
   reg _399916_399916 ; 
   reg __399916_399916;
   reg _399917_399917 ; 
   reg __399917_399917;
   reg _399918_399918 ; 
   reg __399918_399918;
   reg _399919_399919 ; 
   reg __399919_399919;
   reg _399920_399920 ; 
   reg __399920_399920;
   reg _399921_399921 ; 
   reg __399921_399921;
   reg _399922_399922 ; 
   reg __399922_399922;
   reg _399923_399923 ; 
   reg __399923_399923;
   reg _399924_399924 ; 
   reg __399924_399924;
   reg _399925_399925 ; 
   reg __399925_399925;
   reg _399926_399926 ; 
   reg __399926_399926;
   reg _399927_399927 ; 
   reg __399927_399927;
   reg _399928_399928 ; 
   reg __399928_399928;
   reg _399929_399929 ; 
   reg __399929_399929;
   reg _399930_399930 ; 
   reg __399930_399930;
   reg _399931_399931 ; 
   reg __399931_399931;
   reg _399932_399932 ; 
   reg __399932_399932;
   reg _399933_399933 ; 
   reg __399933_399933;
   reg _399934_399934 ; 
   reg __399934_399934;
   reg _399935_399935 ; 
   reg __399935_399935;
   reg _399936_399936 ; 
   reg __399936_399936;
   reg _399937_399937 ; 
   reg __399937_399937;
   reg _399938_399938 ; 
   reg __399938_399938;
   reg _399939_399939 ; 
   reg __399939_399939;
   reg _399940_399940 ; 
   reg __399940_399940;
   reg _399941_399941 ; 
   reg __399941_399941;
   reg _399942_399942 ; 
   reg __399942_399942;
   reg _399943_399943 ; 
   reg __399943_399943;
   reg _399944_399944 ; 
   reg __399944_399944;
   reg _399945_399945 ; 
   reg __399945_399945;
   reg _399946_399946 ; 
   reg __399946_399946;
   reg _399947_399947 ; 
   reg __399947_399947;
   reg _399948_399948 ; 
   reg __399948_399948;
   reg _399949_399949 ; 
   reg __399949_399949;
   reg _399950_399950 ; 
   reg __399950_399950;
   reg _399951_399951 ; 
   reg __399951_399951;
   reg _399952_399952 ; 
   reg __399952_399952;
   reg _399953_399953 ; 
   reg __399953_399953;
   reg _399954_399954 ; 
   reg __399954_399954;
   reg _399955_399955 ; 
   reg __399955_399955;
   reg _399956_399956 ; 
   reg __399956_399956;
   reg _399957_399957 ; 
   reg __399957_399957;
   reg _399958_399958 ; 
   reg __399958_399958;
   reg _399959_399959 ; 
   reg __399959_399959;
   reg _399960_399960 ; 
   reg __399960_399960;
   reg _399961_399961 ; 
   reg __399961_399961;
   reg _399962_399962 ; 
   reg __399962_399962;
   reg _399963_399963 ; 
   reg __399963_399963;
   reg _399964_399964 ; 
   reg __399964_399964;
   reg _399965_399965 ; 
   reg __399965_399965;
   reg _399966_399966 ; 
   reg __399966_399966;
   reg _399967_399967 ; 
   reg __399967_399967;
   reg _399968_399968 ; 
   reg __399968_399968;
   reg _399969_399969 ; 
   reg __399969_399969;
   reg _399970_399970 ; 
   reg __399970_399970;
   reg _399971_399971 ; 
   reg __399971_399971;
   reg _399972_399972 ; 
   reg __399972_399972;
   reg _399973_399973 ; 
   reg __399973_399973;
   reg _399974_399974 ; 
   reg __399974_399974;
   reg _399975_399975 ; 
   reg __399975_399975;
   reg _399976_399976 ; 
   reg __399976_399976;
   reg _399977_399977 ; 
   reg __399977_399977;
   reg _399978_399978 ; 
   reg __399978_399978;
   reg _399979_399979 ; 
   reg __399979_399979;
   reg _399980_399980 ; 
   reg __399980_399980;
   reg _399981_399981 ; 
   reg __399981_399981;
   reg _399982_399982 ; 
   reg __399982_399982;
   reg _399983_399983 ; 
   reg __399983_399983;
   reg _399984_399984 ; 
   reg __399984_399984;
   reg _399985_399985 ; 
   reg __399985_399985;
   reg _399986_399986 ; 
   reg __399986_399986;
   reg _399987_399987 ; 
   reg __399987_399987;
   reg _399988_399988 ; 
   reg __399988_399988;
   reg _399989_399989 ; 
   reg __399989_399989;
   reg _399990_399990 ; 
   reg __399990_399990;
   reg _399991_399991 ; 
   reg __399991_399991;
   reg _399992_399992 ; 
   reg __399992_399992;
   reg _399993_399993 ; 
   reg __399993_399993;
   reg _399994_399994 ; 
   reg __399994_399994;
   reg _399995_399995 ; 
   reg __399995_399995;
   reg _399996_399996 ; 
   reg __399996_399996;
   reg _399997_399997 ; 
   reg __399997_399997;
   reg _399998_399998 ; 
   reg __399998_399998;
   reg _399999_399999 ; 
   reg __399999_399999;
   reg _400000_400000 ; 
   reg __400000_400000;
   reg _400001_400001 ; 
   reg __400001_400001;
   reg _400002_400002 ; 
   reg __400002_400002;
   reg _400003_400003 ; 
   reg __400003_400003;
   reg _400004_400004 ; 
   reg __400004_400004;
   reg _400005_400005 ; 
   reg __400005_400005;
   reg _400006_400006 ; 
   reg __400006_400006;
   reg _400007_400007 ; 
   reg __400007_400007;
   reg _400008_400008 ; 
   reg __400008_400008;
   reg _400009_400009 ; 
   reg __400009_400009;
   reg _400010_400010 ; 
   reg __400010_400010;
   reg _400011_400011 ; 
   reg __400011_400011;
   reg _400012_400012 ; 
   reg __400012_400012;
   reg _400013_400013 ; 
   reg __400013_400013;
   reg _400014_400014 ; 
   reg __400014_400014;
   reg _400015_400015 ; 
   reg __400015_400015;
   reg _400016_400016 ; 
   reg __400016_400016;
   reg _400017_400017 ; 
   reg __400017_400017;
   reg _400018_400018 ; 
   reg __400018_400018;
   reg _400019_400019 ; 
   reg __400019_400019;
   reg _400020_400020 ; 
   reg __400020_400020;
   reg _400021_400021 ; 
   reg __400021_400021;
   reg _400022_400022 ; 
   reg __400022_400022;
   reg _400023_400023 ; 
   reg __400023_400023;
   reg _400024_400024 ; 
   reg __400024_400024;
   reg _400025_400025 ; 
   reg __400025_400025;
   reg _400026_400026 ; 
   reg __400026_400026;
   reg _400027_400027 ; 
   reg __400027_400027;
   reg _400028_400028 ; 
   reg __400028_400028;
   reg _400029_400029 ; 
   reg __400029_400029;
   reg _400030_400030 ; 
   reg __400030_400030;
   reg _400031_400031 ; 
   reg __400031_400031;
   reg _400032_400032 ; 
   reg __400032_400032;
   reg _400033_400033 ; 
   reg __400033_400033;
   reg _400034_400034 ; 
   reg __400034_400034;
   reg _400035_400035 ; 
   reg __400035_400035;
   reg _400036_400036 ; 
   reg __400036_400036;
   reg _400037_400037 ; 
   reg __400037_400037;
   reg _400038_400038 ; 
   reg __400038_400038;
   reg _400039_400039 ; 
   reg __400039_400039;
   reg _400040_400040 ; 
   reg __400040_400040;
   reg _400041_400041 ; 
   reg __400041_400041;
   reg _400042_400042 ; 
   reg __400042_400042;
   reg _400043_400043 ; 
   reg __400043_400043;
   reg _400044_400044 ; 
   reg __400044_400044;
   reg _400045_400045 ; 
   reg __400045_400045;
   reg _400046_400046 ; 
   reg __400046_400046;
   reg _400047_400047 ; 
   reg __400047_400047;
   reg _400048_400048 ; 
   reg __400048_400048;
   reg _400049_400049 ; 
   reg __400049_400049;
   reg _400050_400050 ; 
   reg __400050_400050;
   reg _400051_400051 ; 
   reg __400051_400051;
   reg _400052_400052 ; 
   reg __400052_400052;
   reg _400053_400053 ; 
   reg __400053_400053;
   reg _400054_400054 ; 
   reg __400054_400054;
   reg _400055_400055 ; 
   reg __400055_400055;
   reg _400056_400056 ; 
   reg __400056_400056;
   reg _400057_400057 ; 
   reg __400057_400057;
   reg _400058_400058 ; 
   reg __400058_400058;
   reg _400059_400059 ; 
   reg __400059_400059;
   reg _400060_400060 ; 
   reg __400060_400060;
   reg _400061_400061 ; 
   reg __400061_400061;
   reg _400062_400062 ; 
   reg __400062_400062;
   reg _400063_400063 ; 
   reg __400063_400063;
   reg _400064_400064 ; 
   reg __400064_400064;
   reg _400065_400065 ; 
   reg __400065_400065;
   reg _400066_400066 ; 
   reg __400066_400066;
   reg _400067_400067 ; 
   reg __400067_400067;
   reg _400068_400068 ; 
   reg __400068_400068;
   reg _400069_400069 ; 
   reg __400069_400069;
   reg _400070_400070 ; 
   reg __400070_400070;
   reg _400071_400071 ; 
   reg __400071_400071;
   reg _400072_400072 ; 
   reg __400072_400072;
   reg _400073_400073 ; 
   reg __400073_400073;
   reg _400074_400074 ; 
   reg __400074_400074;
   reg _400075_400075 ; 
   reg __400075_400075;
   reg _400076_400076 ; 
   reg __400076_400076;
   reg _400077_400077 ; 
   reg __400077_400077;
   reg _400078_400078 ; 
   reg __400078_400078;
   reg _400079_400079 ; 
   reg __400079_400079;
   reg _400080_400080 ; 
   reg __400080_400080;
   reg _400081_400081 ; 
   reg __400081_400081;
   reg _400082_400082 ; 
   reg __400082_400082;
   reg _400083_400083 ; 
   reg __400083_400083;
   reg _400084_400084 ; 
   reg __400084_400084;
   reg _400085_400085 ; 
   reg __400085_400085;
   reg _400086_400086 ; 
   reg __400086_400086;
   reg _400087_400087 ; 
   reg __400087_400087;
   reg _400088_400088 ; 
   reg __400088_400088;
   reg _400089_400089 ; 
   reg __400089_400089;
   reg _400090_400090 ; 
   reg __400090_400090;
   reg _400091_400091 ; 
   reg __400091_400091;
   reg _400092_400092 ; 
   reg __400092_400092;
   reg _400093_400093 ; 
   reg __400093_400093;
   reg _400094_400094 ; 
   reg __400094_400094;
   reg _400095_400095 ; 
   reg __400095_400095;
   reg _400096_400096 ; 
   reg __400096_400096;
   reg _400097_400097 ; 
   reg __400097_400097;
   reg _400098_400098 ; 
   reg __400098_400098;
   reg _400099_400099 ; 
   reg __400099_400099;
   reg _400100_400100 ; 
   reg __400100_400100;
   reg _400101_400101 ; 
   reg __400101_400101;
   reg _400102_400102 ; 
   reg __400102_400102;
   reg _400103_400103 ; 
   reg __400103_400103;
   reg _400104_400104 ; 
   reg __400104_400104;
   reg _400105_400105 ; 
   reg __400105_400105;
   reg _400106_400106 ; 
   reg __400106_400106;
   reg _400107_400107 ; 
   reg __400107_400107;
   reg _400108_400108 ; 
   reg __400108_400108;
   reg _400109_400109 ; 
   reg __400109_400109;
   reg _400110_400110 ; 
   reg __400110_400110;
   reg _400111_400111 ; 
   reg __400111_400111;
   reg _400112_400112 ; 
   reg __400112_400112;
   reg _400113_400113 ; 
   reg __400113_400113;
   reg _400114_400114 ; 
   reg __400114_400114;
   reg _400115_400115 ; 
   reg __400115_400115;
   reg _400116_400116 ; 
   reg __400116_400116;
   reg _400117_400117 ; 
   reg __400117_400117;
   reg _400118_400118 ; 
   reg __400118_400118;
   reg _400119_400119 ; 
   reg __400119_400119;
   reg _400120_400120 ; 
   reg __400120_400120;
   reg _400121_400121 ; 
   reg __400121_400121;
   reg _400122_400122 ; 
   reg __400122_400122;
   reg _400123_400123 ; 
   reg __400123_400123;
   reg _400124_400124 ; 
   reg __400124_400124;
   reg _400125_400125 ; 
   reg __400125_400125;
   reg _400126_400126 ; 
   reg __400126_400126;
   reg _400127_400127 ; 
   reg __400127_400127;
   reg _400128_400128 ; 
   reg __400128_400128;
   reg _400129_400129 ; 
   reg __400129_400129;
   reg _400130_400130 ; 
   reg __400130_400130;
   reg _400131_400131 ; 
   reg __400131_400131;
   reg _400132_400132 ; 
   reg __400132_400132;
   reg _400133_400133 ; 
   reg __400133_400133;
   reg _400134_400134 ; 
   reg __400134_400134;
   reg _400135_400135 ; 
   reg __400135_400135;
   reg _400136_400136 ; 
   reg __400136_400136;
   reg _400137_400137 ; 
   reg __400137_400137;
   reg _400138_400138 ; 
   reg __400138_400138;
   reg _400139_400139 ; 
   reg __400139_400139;
   reg _400140_400140 ; 
   reg __400140_400140;
   reg _400141_400141 ; 
   reg __400141_400141;
   reg _400142_400142 ; 
   reg __400142_400142;
   reg _400143_400143 ; 
   reg __400143_400143;
   reg _400144_400144 ; 
   reg __400144_400144;
   reg _400145_400145 ; 
   reg __400145_400145;
   reg _400146_400146 ; 
   reg __400146_400146;
   reg _400147_400147 ; 
   reg __400147_400147;
   reg _400148_400148 ; 
   reg __400148_400148;
   reg _400149_400149 ; 
   reg __400149_400149;
   reg _400150_400150 ; 
   reg __400150_400150;
   reg _400151_400151 ; 
   reg __400151_400151;
   reg _400152_400152 ; 
   reg __400152_400152;
   reg _400153_400153 ; 
   reg __400153_400153;
   reg _400154_400154 ; 
   reg __400154_400154;
   reg _400155_400155 ; 
   reg __400155_400155;
   reg _400156_400156 ; 
   reg __400156_400156;
   reg _400157_400157 ; 
   reg __400157_400157;
   reg _400158_400158 ; 
   reg __400158_400158;
   reg _400159_400159 ; 
   reg __400159_400159;
   reg _400160_400160 ; 
   reg __400160_400160;
   reg _400161_400161 ; 
   reg __400161_400161;
   reg _400162_400162 ; 
   reg __400162_400162;
   reg _400163_400163 ; 
   reg __400163_400163;
   reg _400164_400164 ; 
   reg __400164_400164;
   reg _400165_400165 ; 
   reg __400165_400165;
   reg _400166_400166 ; 
   reg __400166_400166;
   reg _400167_400167 ; 
   reg __400167_400167;
   reg _400168_400168 ; 
   reg __400168_400168;
   reg _400169_400169 ; 
   reg __400169_400169;
   reg _400170_400170 ; 
   reg __400170_400170;
   reg _400171_400171 ; 
   reg __400171_400171;
   reg _400172_400172 ; 
   reg __400172_400172;
   reg _400173_400173 ; 
   reg __400173_400173;
   reg _400174_400174 ; 
   reg __400174_400174;
   reg _400175_400175 ; 
   reg __400175_400175;
   reg _400176_400176 ; 
   reg __400176_400176;
   reg _400177_400177 ; 
   reg __400177_400177;
   reg _400178_400178 ; 
   reg __400178_400178;
   reg _400179_400179 ; 
   reg __400179_400179;
   reg _400180_400180 ; 
   reg __400180_400180;
   reg _400181_400181 ; 
   reg __400181_400181;
   reg _400182_400182 ; 
   reg __400182_400182;
   reg _400183_400183 ; 
   reg __400183_400183;
   reg _400184_400184 ; 
   reg __400184_400184;
   reg _400185_400185 ; 
   reg __400185_400185;
   reg _400186_400186 ; 
   reg __400186_400186;
   reg _400187_400187 ; 
   reg __400187_400187;
   reg _400188_400188 ; 
   reg __400188_400188;
   reg _400189_400189 ; 
   reg __400189_400189;
   reg _400190_400190 ; 
   reg __400190_400190;
   reg _400191_400191 ; 
   reg __400191_400191;
   reg _400192_400192 ; 
   reg __400192_400192;
   reg _400193_400193 ; 
   reg __400193_400193;
   reg _400194_400194 ; 
   reg __400194_400194;
   reg _400195_400195 ; 
   reg __400195_400195;
   reg _400196_400196 ; 
   reg __400196_400196;
   reg _400197_400197 ; 
   reg __400197_400197;
   reg _400198_400198 ; 
   reg __400198_400198;
   reg _400199_400199 ; 
   reg __400199_400199;
   reg _400200_400200 ; 
   reg __400200_400200;
   reg _400201_400201 ; 
   reg __400201_400201;
   reg _400202_400202 ; 
   reg __400202_400202;
   reg _400203_400203 ; 
   reg __400203_400203;
   reg _400204_400204 ; 
   reg __400204_400204;
   reg _400205_400205 ; 
   reg __400205_400205;
   reg _400206_400206 ; 
   reg __400206_400206;
   reg _400207_400207 ; 
   reg __400207_400207;
   reg _400208_400208 ; 
   reg __400208_400208;
   reg _400209_400209 ; 
   reg __400209_400209;
   reg _400210_400210 ; 
   reg __400210_400210;
   reg _400211_400211 ; 
   reg __400211_400211;
   reg _400212_400212 ; 
   reg __400212_400212;
   reg _400213_400213 ; 
   reg __400213_400213;
   reg _400214_400214 ; 
   reg __400214_400214;
   reg _400215_400215 ; 
   reg __400215_400215;
   reg _400216_400216 ; 
   reg __400216_400216;
   reg _400217_400217 ; 
   reg __400217_400217;
   reg _400218_400218 ; 
   reg __400218_400218;
   reg _400219_400219 ; 
   reg __400219_400219;
   reg _400220_400220 ; 
   reg __400220_400220;
   reg _400221_400221 ; 
   reg __400221_400221;
   reg _400222_400222 ; 
   reg __400222_400222;
   reg _400223_400223 ; 
   reg __400223_400223;
   reg _400224_400224 ; 
   reg __400224_400224;
   reg _400225_400225 ; 
   reg __400225_400225;
   reg _400226_400226 ; 
   reg __400226_400226;
   reg _400227_400227 ; 
   reg __400227_400227;
   reg _400228_400228 ; 
   reg __400228_400228;
   reg _400229_400229 ; 
   reg __400229_400229;
   reg _400230_400230 ; 
   reg __400230_400230;
   reg _400231_400231 ; 
   reg __400231_400231;
   reg _400232_400232 ; 
   reg __400232_400232;
   reg _400233_400233 ; 
   reg __400233_400233;
   reg _400234_400234 ; 
   reg __400234_400234;
   reg _400235_400235 ; 
   reg __400235_400235;
   reg _400236_400236 ; 
   reg __400236_400236;
   reg _400237_400237 ; 
   reg __400237_400237;
   reg _400238_400238 ; 
   reg __400238_400238;
   reg _400239_400239 ; 
   reg __400239_400239;
   reg _400240_400240 ; 
   reg __400240_400240;
   reg _400241_400241 ; 
   reg __400241_400241;
   reg _400242_400242 ; 
   reg __400242_400242;
   reg _400243_400243 ; 
   reg __400243_400243;
   reg _400244_400244 ; 
   reg __400244_400244;
   reg _400245_400245 ; 
   reg __400245_400245;
   reg _400246_400246 ; 
   reg __400246_400246;
   reg _400247_400247 ; 
   reg __400247_400247;
   reg _400248_400248 ; 
   reg __400248_400248;
   reg _400249_400249 ; 
   reg __400249_400249;
   reg _400250_400250 ; 
   reg __400250_400250;
   reg _400251_400251 ; 
   reg __400251_400251;
   reg _400252_400252 ; 
   reg __400252_400252;
   reg _400253_400253 ; 
   reg __400253_400253;
   reg _400254_400254 ; 
   reg __400254_400254;
   reg _400255_400255 ; 
   reg __400255_400255;
   reg _400256_400256 ; 
   reg __400256_400256;
   reg _400257_400257 ; 
   reg __400257_400257;
   reg _400258_400258 ; 
   reg __400258_400258;
   reg _400259_400259 ; 
   reg __400259_400259;
   reg _400260_400260 ; 
   reg __400260_400260;
   reg _400261_400261 ; 
   reg __400261_400261;
   reg _400262_400262 ; 
   reg __400262_400262;
   reg _400263_400263 ; 
   reg __400263_400263;
   reg _400264_400264 ; 
   reg __400264_400264;
   reg _400265_400265 ; 
   reg __400265_400265;
   reg _400266_400266 ; 
   reg __400266_400266;
   reg _400267_400267 ; 
   reg __400267_400267;
   reg _400268_400268 ; 
   reg __400268_400268;
   reg _400269_400269 ; 
   reg __400269_400269;
   reg _400270_400270 ; 
   reg __400270_400270;
   reg _400271_400271 ; 
   reg __400271_400271;
   reg _400272_400272 ; 
   reg __400272_400272;
   reg _400273_400273 ; 
   reg __400273_400273;
   reg _400274_400274 ; 
   reg __400274_400274;
   reg _400275_400275 ; 
   reg __400275_400275;
   reg _400276_400276 ; 
   reg __400276_400276;
   reg _400277_400277 ; 
   reg __400277_400277;
   reg _400278_400278 ; 
   reg __400278_400278;
   reg _400279_400279 ; 
   reg __400279_400279;
   reg _400280_400280 ; 
   reg __400280_400280;
   reg _400281_400281 ; 
   reg __400281_400281;
   reg _400282_400282 ; 
   reg __400282_400282;
   reg _400283_400283 ; 
   reg __400283_400283;
   reg _400284_400284 ; 
   reg __400284_400284;
   reg _400285_400285 ; 
   reg __400285_400285;
   reg _400286_400286 ; 
   reg __400286_400286;
   reg _400287_400287 ; 
   reg __400287_400287;
   reg _400288_400288 ; 
   reg __400288_400288;
   reg _400289_400289 ; 
   reg __400289_400289;
   reg _400290_400290 ; 
   reg __400290_400290;
   reg _400291_400291 ; 
   reg __400291_400291;
   reg _400292_400292 ; 
   reg __400292_400292;
   reg _400293_400293 ; 
   reg __400293_400293;
   reg _400294_400294 ; 
   reg __400294_400294;
   reg _400295_400295 ; 
   reg __400295_400295;
   reg _400296_400296 ; 
   reg __400296_400296;
   reg _400297_400297 ; 
   reg __400297_400297;
   reg _400298_400298 ; 
   reg __400298_400298;
   reg _400299_400299 ; 
   reg __400299_400299;
   reg _400300_400300 ; 
   reg __400300_400300;
   reg _400301_400301 ; 
   reg __400301_400301;
   reg _400302_400302 ; 
   reg __400302_400302;
   reg _400303_400303 ; 
   reg __400303_400303;
   reg _400304_400304 ; 
   reg __400304_400304;
   reg _400305_400305 ; 
   reg __400305_400305;
   reg _400306_400306 ; 
   reg __400306_400306;
   reg _400307_400307 ; 
   reg __400307_400307;
   reg _400308_400308 ; 
   reg __400308_400308;
   reg _400309_400309 ; 
   reg __400309_400309;
   reg _400310_400310 ; 
   reg __400310_400310;
   reg _400311_400311 ; 
   reg __400311_400311;
   reg _400312_400312 ; 
   reg __400312_400312;
   reg _400313_400313 ; 
   reg __400313_400313;
   reg _400314_400314 ; 
   reg __400314_400314;
   reg _400315_400315 ; 
   reg __400315_400315;
   reg _400316_400316 ; 
   reg __400316_400316;
   reg _400317_400317 ; 
   reg __400317_400317;
   reg _400318_400318 ; 
   reg __400318_400318;
   reg _400319_400319 ; 
   reg __400319_400319;
   reg _400320_400320 ; 
   reg __400320_400320;
   reg _400321_400321 ; 
   reg __400321_400321;
   reg _400322_400322 ; 
   reg __400322_400322;
   reg _400323_400323 ; 
   reg __400323_400323;
   reg _400324_400324 ; 
   reg __400324_400324;
   reg _400325_400325 ; 
   reg __400325_400325;
   reg _400326_400326 ; 
   reg __400326_400326;
   reg _400327_400327 ; 
   reg __400327_400327;
   reg _400328_400328 ; 
   reg __400328_400328;
   reg _400329_400329 ; 
   reg __400329_400329;
   reg _400330_400330 ; 
   reg __400330_400330;
   reg _400331_400331 ; 
   reg __400331_400331;
   reg _400332_400332 ; 
   reg __400332_400332;
   reg _400333_400333 ; 
   reg __400333_400333;
   reg _400334_400334 ; 
   reg __400334_400334;
   reg _400335_400335 ; 
   reg __400335_400335;
   reg _400336_400336 ; 
   reg __400336_400336;
   reg _400337_400337 ; 
   reg __400337_400337;
   reg _400338_400338 ; 
   reg __400338_400338;
   reg _400339_400339 ; 
   reg __400339_400339;
   reg _400340_400340 ; 
   reg __400340_400340;
   reg _400341_400341 ; 
   reg __400341_400341;
   reg _400342_400342 ; 
   reg __400342_400342;
   reg _400343_400343 ; 
   reg __400343_400343;
   reg _400344_400344 ; 
   reg __400344_400344;
   reg _400345_400345 ; 
   reg __400345_400345;
   reg _400346_400346 ; 
   reg __400346_400346;
   reg _400347_400347 ; 
   reg __400347_400347;
   reg _400348_400348 ; 
   reg __400348_400348;
   reg _400349_400349 ; 
   reg __400349_400349;
   reg _400350_400350 ; 
   reg __400350_400350;
   reg _400351_400351 ; 
   reg __400351_400351;
   reg _400352_400352 ; 
   reg __400352_400352;
   reg _400353_400353 ; 
   reg __400353_400353;
   reg _400354_400354 ; 
   reg __400354_400354;
   reg _400355_400355 ; 
   reg __400355_400355;
   reg _400356_400356 ; 
   reg __400356_400356;
   reg _400357_400357 ; 
   reg __400357_400357;
   reg _400358_400358 ; 
   reg __400358_400358;
   reg _400359_400359 ; 
   reg __400359_400359;
   reg _400360_400360 ; 
   reg __400360_400360;
   reg _400361_400361 ; 
   reg __400361_400361;
   reg _400362_400362 ; 
   reg __400362_400362;
   reg _400363_400363 ; 
   reg __400363_400363;
   reg _400364_400364 ; 
   reg __400364_400364;
   reg _400365_400365 ; 
   reg __400365_400365;
   reg _400366_400366 ; 
   reg __400366_400366;
   reg _400367_400367 ; 
   reg __400367_400367;
   reg _400368_400368 ; 
   reg __400368_400368;
   reg _400369_400369 ; 
   reg __400369_400369;
   reg _400370_400370 ; 
   reg __400370_400370;
   reg _400371_400371 ; 
   reg __400371_400371;
   reg _400372_400372 ; 
   reg __400372_400372;
   reg _400373_400373 ; 
   reg __400373_400373;
   reg _400374_400374 ; 
   reg __400374_400374;
   reg _400375_400375 ; 
   reg __400375_400375;
   reg _400376_400376 ; 
   reg __400376_400376;
   reg _400377_400377 ; 
   reg __400377_400377;
   reg _400378_400378 ; 
   reg __400378_400378;
   reg _400379_400379 ; 
   reg __400379_400379;
   reg _400380_400380 ; 
   reg __400380_400380;
   reg _400381_400381 ; 
   reg __400381_400381;
   reg _400382_400382 ; 
   reg __400382_400382;
   reg _400383_400383 ; 
   reg __400383_400383;
   reg _400384_400384 ; 
   reg __400384_400384;
   reg _400385_400385 ; 
   reg __400385_400385;
   reg _400386_400386 ; 
   reg __400386_400386;
   reg _400387_400387 ; 
   reg __400387_400387;
   reg _400388_400388 ; 
   reg __400388_400388;
   reg _400389_400389 ; 
   reg __400389_400389;
   reg _400390_400390 ; 
   reg __400390_400390;
   reg _400391_400391 ; 
   reg __400391_400391;
   reg _400392_400392 ; 
   reg __400392_400392;
   reg _400393_400393 ; 
   reg __400393_400393;
   reg _400394_400394 ; 
   reg __400394_400394;
   reg _400395_400395 ; 
   reg __400395_400395;
   reg _400396_400396 ; 
   reg __400396_400396;
   reg _400397_400397 ; 
   reg __400397_400397;
   reg _400398_400398 ; 
   reg __400398_400398;
   reg _400399_400399 ; 
   reg __400399_400399;
   reg _400400_400400 ; 
   reg __400400_400400;
   reg _400401_400401 ; 
   reg __400401_400401;
   reg _400402_400402 ; 
   reg __400402_400402;
   reg _400403_400403 ; 
   reg __400403_400403;
   reg _400404_400404 ; 
   reg __400404_400404;
   reg _400405_400405 ; 
   reg __400405_400405;
   reg _400406_400406 ; 
   reg __400406_400406;
   reg _400407_400407 ; 
   reg __400407_400407;
   reg _400408_400408 ; 
   reg __400408_400408;
   reg _400409_400409 ; 
   reg __400409_400409;
   reg _400410_400410 ; 
   reg __400410_400410;
   reg _400411_400411 ; 
   reg __400411_400411;
   reg _400412_400412 ; 
   reg __400412_400412;
   reg _400413_400413 ; 
   reg __400413_400413;
   reg _400414_400414 ; 
   reg __400414_400414;
   reg _400415_400415 ; 
   reg __400415_400415;
   reg _400416_400416 ; 
   reg __400416_400416;
   reg _400417_400417 ; 
   reg __400417_400417;
   reg _400418_400418 ; 
   reg __400418_400418;
   reg _400419_400419 ; 
   reg __400419_400419;
   reg _400420_400420 ; 
   reg __400420_400420;
   reg _400421_400421 ; 
   reg __400421_400421;
   reg _400422_400422 ; 
   reg __400422_400422;
   reg _400423_400423 ; 
   reg __400423_400423;
   reg _400424_400424 ; 
   reg __400424_400424;
   reg _400425_400425 ; 
   reg __400425_400425;
   reg _400426_400426 ; 
   reg __400426_400426;
   reg _400427_400427 ; 
   reg __400427_400427;
   reg _400428_400428 ; 
   reg __400428_400428;
   reg _400429_400429 ; 
   reg __400429_400429;
   reg _400430_400430 ; 
   reg __400430_400430;
   reg _400431_400431 ; 
   reg __400431_400431;
   reg _400432_400432 ; 
   reg __400432_400432;
   reg _400433_400433 ; 
   reg __400433_400433;
   reg _400434_400434 ; 
   reg __400434_400434;
   reg _400435_400435 ; 
   reg __400435_400435;
   reg _400436_400436 ; 
   reg __400436_400436;
   reg _400437_400437 ; 
   reg __400437_400437;
   reg _400438_400438 ; 
   reg __400438_400438;
   reg _400439_400439 ; 
   reg __400439_400439;
   reg _400440_400440 ; 
   reg __400440_400440;
   reg _400441_400441 ; 
   reg __400441_400441;
   reg _400442_400442 ; 
   reg __400442_400442;
   reg _400443_400443 ; 
   reg __400443_400443;
   reg _400444_400444 ; 
   reg __400444_400444;
   reg _400445_400445 ; 
   reg __400445_400445;
   reg _400446_400446 ; 
   reg __400446_400446;
   reg _400447_400447 ; 
   reg __400447_400447;
   reg _400448_400448 ; 
   reg __400448_400448;
   reg _400449_400449 ; 
   reg __400449_400449;
   reg _400450_400450 ; 
   reg __400450_400450;
   reg _400451_400451 ; 
   reg __400451_400451;
   reg _400452_400452 ; 
   reg __400452_400452;
   reg _400453_400453 ; 
   reg __400453_400453;
   reg _400454_400454 ; 
   reg __400454_400454;
   reg _400455_400455 ; 
   reg __400455_400455;
   reg _400456_400456 ; 
   reg __400456_400456;
   reg _400457_400457 ; 
   reg __400457_400457;
   reg _400458_400458 ; 
   reg __400458_400458;
   reg _400459_400459 ; 
   reg __400459_400459;
   reg _400460_400460 ; 
   reg __400460_400460;
   reg _400461_400461 ; 
   reg __400461_400461;
   reg _400462_400462 ; 
   reg __400462_400462;
   reg _400463_400463 ; 
   reg __400463_400463;
   reg _400464_400464 ; 
   reg __400464_400464;
   reg _400465_400465 ; 
   reg __400465_400465;
   reg _400466_400466 ; 
   reg __400466_400466;
   reg _400467_400467 ; 
   reg __400467_400467;
   reg _400468_400468 ; 
   reg __400468_400468;
   reg _400469_400469 ; 
   reg __400469_400469;
   reg _400470_400470 ; 
   reg __400470_400470;
   reg _400471_400471 ; 
   reg __400471_400471;
   reg _400472_400472 ; 
   reg __400472_400472;
   reg _400473_400473 ; 
   reg __400473_400473;
   reg _400474_400474 ; 
   reg __400474_400474;
   reg _400475_400475 ; 
   reg __400475_400475;
   reg _400476_400476 ; 
   reg __400476_400476;
   reg _400477_400477 ; 
   reg __400477_400477;
   reg _400478_400478 ; 
   reg __400478_400478;
   reg _400479_400479 ; 
   reg __400479_400479;
   reg _400480_400480 ; 
   reg __400480_400480;
   reg _400481_400481 ; 
   reg __400481_400481;
   reg _400482_400482 ; 
   reg __400482_400482;
   reg _400483_400483 ; 
   reg __400483_400483;
   reg _400484_400484 ; 
   reg __400484_400484;
   reg _400485_400485 ; 
   reg __400485_400485;
   reg _400486_400486 ; 
   reg __400486_400486;
   reg _400487_400487 ; 
   reg __400487_400487;
   reg _400488_400488 ; 
   reg __400488_400488;
   reg _400489_400489 ; 
   reg __400489_400489;
   reg _400490_400490 ; 
   reg __400490_400490;
   reg _400491_400491 ; 
   reg __400491_400491;
   reg _400492_400492 ; 
   reg __400492_400492;
   reg _400493_400493 ; 
   reg __400493_400493;
   reg _400494_400494 ; 
   reg __400494_400494;
   reg _400495_400495 ; 
   reg __400495_400495;
   reg _400496_400496 ; 
   reg __400496_400496;
   reg _400497_400497 ; 
   reg __400497_400497;
   reg _400498_400498 ; 
   reg __400498_400498;
   reg _400499_400499 ; 
   reg __400499_400499;
   reg _400500_400500 ; 
   reg __400500_400500;
   reg _400501_400501 ; 
   reg __400501_400501;
   reg _400502_400502 ; 
   reg __400502_400502;
   reg _400503_400503 ; 
   reg __400503_400503;
   reg _400504_400504 ; 
   reg __400504_400504;
   reg _400505_400505 ; 
   reg __400505_400505;
   reg _400506_400506 ; 
   reg __400506_400506;
   reg _400507_400507 ; 
   reg __400507_400507;
   reg _400508_400508 ; 
   reg __400508_400508;
   reg _400509_400509 ; 
   reg __400509_400509;
   reg _400510_400510 ; 
   reg __400510_400510;
   reg _400511_400511 ; 
   reg __400511_400511;
   reg _400512_400512 ; 
   reg __400512_400512;
   reg _400513_400513 ; 
   reg __400513_400513;
   reg _400514_400514 ; 
   reg __400514_400514;
   reg _400515_400515 ; 
   reg __400515_400515;
   reg _400516_400516 ; 
   reg __400516_400516;
   reg _400517_400517 ; 
   reg __400517_400517;
   reg _400518_400518 ; 
   reg __400518_400518;
   reg _400519_400519 ; 
   reg __400519_400519;
   reg _400520_400520 ; 
   reg __400520_400520;
   reg _400521_400521 ; 
   reg __400521_400521;
   reg _400522_400522 ; 
   reg __400522_400522;
   reg _400523_400523 ; 
   reg __400523_400523;
   reg _400524_400524 ; 
   reg __400524_400524;
   reg _400525_400525 ; 
   reg __400525_400525;
   reg _400526_400526 ; 
   reg __400526_400526;
   reg _400527_400527 ; 
   reg __400527_400527;
   reg _400528_400528 ; 
   reg __400528_400528;
   reg _400529_400529 ; 
   reg __400529_400529;
   reg _400530_400530 ; 
   reg __400530_400530;
   reg _400531_400531 ; 
   reg __400531_400531;
   reg _400532_400532 ; 
   reg __400532_400532;
   reg _400533_400533 ; 
   reg __400533_400533;
   reg _400534_400534 ; 
   reg __400534_400534;
   reg _400535_400535 ; 
   reg __400535_400535;
   reg _400536_400536 ; 
   reg __400536_400536;
   reg _400537_400537 ; 
   reg __400537_400537;
   reg _400538_400538 ; 
   reg __400538_400538;
   reg _400539_400539 ; 
   reg __400539_400539;
   reg _400540_400540 ; 
   reg __400540_400540;
   reg _400541_400541 ; 
   reg __400541_400541;
   reg _400542_400542 ; 
   reg __400542_400542;
   reg _400543_400543 ; 
   reg __400543_400543;
   reg _400544_400544 ; 
   reg __400544_400544;
   reg _400545_400545 ; 
   reg __400545_400545;
   reg _400546_400546 ; 
   reg __400546_400546;
   reg _400547_400547 ; 
   reg __400547_400547;
   reg _400548_400548 ; 
   reg __400548_400548;
   reg _400549_400549 ; 
   reg __400549_400549;
   reg _400550_400550 ; 
   reg __400550_400550;
   reg _400551_400551 ; 
   reg __400551_400551;
   reg _400552_400552 ; 
   reg __400552_400552;
   reg _400553_400553 ; 
   reg __400553_400553;
   reg _400554_400554 ; 
   reg __400554_400554;
   reg _400555_400555 ; 
   reg __400555_400555;
   reg _400556_400556 ; 
   reg __400556_400556;
   reg _400557_400557 ; 
   reg __400557_400557;
   reg _400558_400558 ; 
   reg __400558_400558;
   reg _400559_400559 ; 
   reg __400559_400559;
   reg _400560_400560 ; 
   reg __400560_400560;
   reg _400561_400561 ; 
   reg __400561_400561;
   reg _400562_400562 ; 
   reg __400562_400562;
   reg _400563_400563 ; 
   reg __400563_400563;
   reg _400564_400564 ; 
   reg __400564_400564;
   reg _400565_400565 ; 
   reg __400565_400565;
   reg _400566_400566 ; 
   reg __400566_400566;
   reg _400567_400567 ; 
   reg __400567_400567;
   reg _400568_400568 ; 
   reg __400568_400568;
   reg _400569_400569 ; 
   reg __400569_400569;
   reg _400570_400570 ; 
   reg __400570_400570;
   reg _400571_400571 ; 
   reg __400571_400571;
   reg _400572_400572 ; 
   reg __400572_400572;
   reg _400573_400573 ; 
   reg __400573_400573;
   reg _400574_400574 ; 
   reg __400574_400574;
   reg _400575_400575 ; 
   reg __400575_400575;
   reg _400576_400576 ; 
   reg __400576_400576;
   reg _400577_400577 ; 
   reg __400577_400577;
   reg _400578_400578 ; 
   reg __400578_400578;
   reg _400579_400579 ; 
   reg __400579_400579;
   reg _400580_400580 ; 
   reg __400580_400580;
   reg _400581_400581 ; 
   reg __400581_400581;
   reg _400582_400582 ; 
   reg __400582_400582;
   reg _400583_400583 ; 
   reg __400583_400583;
   reg _400584_400584 ; 
   reg __400584_400584;
   reg _400585_400585 ; 
   reg __400585_400585;
   reg _400586_400586 ; 
   reg __400586_400586;
   reg _400587_400587 ; 
   reg __400587_400587;
   reg _400588_400588 ; 
   reg __400588_400588;
   reg _400589_400589 ; 
   reg __400589_400589;
   reg _400590_400590 ; 
   reg __400590_400590;
   reg _400591_400591 ; 
   reg __400591_400591;
   reg _400592_400592 ; 
   reg __400592_400592;
   reg _400593_400593 ; 
   reg __400593_400593;
   reg _400594_400594 ; 
   reg __400594_400594;
   reg _400595_400595 ; 
   reg __400595_400595;
   reg _400596_400596 ; 
   reg __400596_400596;
   reg _400597_400597 ; 
   reg __400597_400597;
   reg _400598_400598 ; 
   reg __400598_400598;
   reg _400599_400599 ; 
   reg __400599_400599;
   reg _400600_400600 ; 
   reg __400600_400600;
   reg _400601_400601 ; 
   reg __400601_400601;
   reg _400602_400602 ; 
   reg __400602_400602;
   reg _400603_400603 ; 
   reg __400603_400603;
   reg _400604_400604 ; 
   reg __400604_400604;
   reg _400605_400605 ; 
   reg __400605_400605;
   reg _400606_400606 ; 
   reg __400606_400606;
   reg _400607_400607 ; 
   reg __400607_400607;
   reg _400608_400608 ; 
   reg __400608_400608;
   reg _400609_400609 ; 
   reg __400609_400609;
   reg _400610_400610 ; 
   reg __400610_400610;
   reg _400611_400611 ; 
   reg __400611_400611;
   reg _400612_400612 ; 
   reg __400612_400612;
   reg _400613_400613 ; 
   reg __400613_400613;
   reg _400614_400614 ; 
   reg __400614_400614;
   reg _400615_400615 ; 
   reg __400615_400615;
   reg _400616_400616 ; 
   reg __400616_400616;
   reg _400617_400617 ; 
   reg __400617_400617;
   reg _400618_400618 ; 
   reg __400618_400618;
   reg _400619_400619 ; 
   reg __400619_400619;
   reg _400620_400620 ; 
   reg __400620_400620;
   reg _400621_400621 ; 
   reg __400621_400621;
   reg _400622_400622 ; 
   reg __400622_400622;
   reg _400623_400623 ; 
   reg __400623_400623;
   reg _400624_400624 ; 
   reg __400624_400624;
   reg _400625_400625 ; 
   reg __400625_400625;
   reg _400626_400626 ; 
   reg __400626_400626;
   reg _400627_400627 ; 
   reg __400627_400627;
   reg _400628_400628 ; 
   reg __400628_400628;
   reg _400629_400629 ; 
   reg __400629_400629;
   reg _400630_400630 ; 
   reg __400630_400630;
   reg _400631_400631 ; 
   reg __400631_400631;
   reg _400632_400632 ; 
   reg __400632_400632;
   reg _400633_400633 ; 
   reg __400633_400633;
   reg _400634_400634 ; 
   reg __400634_400634;
   reg _400635_400635 ; 
   reg __400635_400635;
   reg _400636_400636 ; 
   reg __400636_400636;
   reg _400637_400637 ; 
   reg __400637_400637;
   reg _400638_400638 ; 
   reg __400638_400638;
   reg _400639_400639 ; 
   reg __400639_400639;
   reg _400640_400640 ; 
   reg __400640_400640;
   reg _400641_400641 ; 
   reg __400641_400641;
   reg _400642_400642 ; 
   reg __400642_400642;
   reg _400643_400643 ; 
   reg __400643_400643;
   reg _400644_400644 ; 
   reg __400644_400644;
   reg _400645_400645 ; 
   reg __400645_400645;
   reg _400646_400646 ; 
   reg __400646_400646;
   reg _400647_400647 ; 
   reg __400647_400647;
   reg _400648_400648 ; 
   reg __400648_400648;
   reg _400649_400649 ; 
   reg __400649_400649;
   reg _400650_400650 ; 
   reg __400650_400650;
   reg _400651_400651 ; 
   reg __400651_400651;
   reg _400652_400652 ; 
   reg __400652_400652;
   reg _400653_400653 ; 
   reg __400653_400653;
   reg _400654_400654 ; 
   reg __400654_400654;
   reg _400655_400655 ; 
   reg __400655_400655;
   reg _400656_400656 ; 
   reg __400656_400656;
   reg _400657_400657 ; 
   reg __400657_400657;
   reg _400658_400658 ; 
   reg __400658_400658;
   reg _400659_400659 ; 
   reg __400659_400659;
   reg _400660_400660 ; 
   reg __400660_400660;
   reg _400661_400661 ; 
   reg __400661_400661;
   reg _400662_400662 ; 
   reg __400662_400662;
   reg _400663_400663 ; 
   reg __400663_400663;
   reg _400664_400664 ; 
   reg __400664_400664;
   reg _400665_400665 ; 
   reg __400665_400665;
   reg _400666_400666 ; 
   reg __400666_400666;
   reg _400667_400667 ; 
   reg __400667_400667;
   reg _400668_400668 ; 
   reg __400668_400668;
   reg _400669_400669 ; 
   reg __400669_400669;
   reg _400670_400670 ; 
   reg __400670_400670;
   reg _400671_400671 ; 
   reg __400671_400671;
   reg _400672_400672 ; 
   reg __400672_400672;
   reg _400673_400673 ; 
   reg __400673_400673;
   reg _400674_400674 ; 
   reg __400674_400674;
   reg _400675_400675 ; 
   reg __400675_400675;
   reg _400676_400676 ; 
   reg __400676_400676;
   reg _400677_400677 ; 
   reg __400677_400677;
   reg _400678_400678 ; 
   reg __400678_400678;
   reg _400679_400679 ; 
   reg __400679_400679;
   reg _400680_400680 ; 
   reg __400680_400680;
   reg _400681_400681 ; 
   reg __400681_400681;
   reg _400682_400682 ; 
   reg __400682_400682;
   reg _400683_400683 ; 
   reg __400683_400683;
   reg _400684_400684 ; 
   reg __400684_400684;
   reg _400685_400685 ; 
   reg __400685_400685;
   reg _400686_400686 ; 
   reg __400686_400686;
   reg _400687_400687 ; 
   reg __400687_400687;
   reg _400688_400688 ; 
   reg __400688_400688;
   reg _400689_400689 ; 
   reg __400689_400689;
   reg _400690_400690 ; 
   reg __400690_400690;
   reg _400691_400691 ; 
   reg __400691_400691;
   reg _400692_400692 ; 
   reg __400692_400692;
   reg _400693_400693 ; 
   reg __400693_400693;
   reg _400694_400694 ; 
   reg __400694_400694;
   reg _400695_400695 ; 
   reg __400695_400695;
   reg _400696_400696 ; 
   reg __400696_400696;
   reg _400697_400697 ; 
   reg __400697_400697;
   reg _400698_400698 ; 
   reg __400698_400698;
   reg _400699_400699 ; 
   reg __400699_400699;
   reg _400700_400700 ; 
   reg __400700_400700;
   reg _400701_400701 ; 
   reg __400701_400701;
   reg _400702_400702 ; 
   reg __400702_400702;
   reg _400703_400703 ; 
   reg __400703_400703;
   reg _400704_400704 ; 
   reg __400704_400704;
   reg _400705_400705 ; 
   reg __400705_400705;
   reg _400706_400706 ; 
   reg __400706_400706;
   reg _400707_400707 ; 
   reg __400707_400707;
   reg _400708_400708 ; 
   reg __400708_400708;
   reg _400709_400709 ; 
   reg __400709_400709;
   reg _400710_400710 ; 
   reg __400710_400710;
   reg _400711_400711 ; 
   reg __400711_400711;
   reg _400712_400712 ; 
   reg __400712_400712;
   reg _400713_400713 ; 
   reg __400713_400713;
   reg _400714_400714 ; 
   reg __400714_400714;
   reg _400715_400715 ; 
   reg __400715_400715;
   reg _400716_400716 ; 
   reg __400716_400716;
   reg _400717_400717 ; 
   reg __400717_400717;
   reg _400718_400718 ; 
   reg __400718_400718;
   reg _400719_400719 ; 
   reg __400719_400719;
   reg _400720_400720 ; 
   reg __400720_400720;
   reg _400721_400721 ; 
   reg __400721_400721;
   reg _400722_400722 ; 
   reg __400722_400722;
   reg _400723_400723 ; 
   reg __400723_400723;
   reg _400724_400724 ; 
   reg __400724_400724;
   reg _400725_400725 ; 
   reg __400725_400725;
   reg _400726_400726 ; 
   reg __400726_400726;
   reg _400727_400727 ; 
   reg __400727_400727;
   reg _400728_400728 ; 
   reg __400728_400728;
   reg _400729_400729 ; 
   reg __400729_400729;
   reg _400730_400730 ; 
   reg __400730_400730;
   reg _400731_400731 ; 
   reg __400731_400731;
   reg _400732_400732 ; 
   reg __400732_400732;
   reg _400733_400733 ; 
   reg __400733_400733;
   reg _400734_400734 ; 
   reg __400734_400734;
   reg _400735_400735 ; 
   reg __400735_400735;
   reg _400736_400736 ; 
   reg __400736_400736;
   reg _400737_400737 ; 
   reg __400737_400737;
   reg _400738_400738 ; 
   reg __400738_400738;
   reg _400739_400739 ; 
   reg __400739_400739;
   reg _400740_400740 ; 
   reg __400740_400740;
   reg _400741_400741 ; 
   reg __400741_400741;
   reg _400742_400742 ; 
   reg __400742_400742;
   reg _400743_400743 ; 
   reg __400743_400743;
   reg _400744_400744 ; 
   reg __400744_400744;
   reg _400745_400745 ; 
   reg __400745_400745;
   reg _400746_400746 ; 
   reg __400746_400746;
   reg _400747_400747 ; 
   reg __400747_400747;
   reg _400748_400748 ; 
   reg __400748_400748;
   reg _400749_400749 ; 
   reg __400749_400749;
   reg _400750_400750 ; 
   reg __400750_400750;
   reg _400751_400751 ; 
   reg __400751_400751;
   reg _400752_400752 ; 
   reg __400752_400752;
   reg _400753_400753 ; 
   reg __400753_400753;
   reg _400754_400754 ; 
   reg __400754_400754;
   reg _400755_400755 ; 
   reg __400755_400755;
   reg _400756_400756 ; 
   reg __400756_400756;
   reg _400757_400757 ; 
   reg __400757_400757;
   reg _400758_400758 ; 
   reg __400758_400758;
   reg _400759_400759 ; 
   reg __400759_400759;
   reg _400760_400760 ; 
   reg __400760_400760;
   reg _400761_400761 ; 
   reg __400761_400761;
   reg _400762_400762 ; 
   reg __400762_400762;
   reg _400763_400763 ; 
   reg __400763_400763;
   reg _400764_400764 ; 
   reg __400764_400764;
   reg _400765_400765 ; 
   reg __400765_400765;
   reg _400766_400766 ; 
   reg __400766_400766;
   reg _400767_400767 ; 
   reg __400767_400767;
   reg _400768_400768 ; 
   reg __400768_400768;
   reg _400769_400769 ; 
   reg __400769_400769;
   reg _400770_400770 ; 
   reg __400770_400770;
   reg _400771_400771 ; 
   reg __400771_400771;
   reg _400772_400772 ; 
   reg __400772_400772;
   reg _400773_400773 ; 
   reg __400773_400773;
   reg _400774_400774 ; 
   reg __400774_400774;
   reg _400775_400775 ; 
   reg __400775_400775;
   reg _400776_400776 ; 
   reg __400776_400776;
   reg _400777_400777 ; 
   reg __400777_400777;
   reg _400778_400778 ; 
   reg __400778_400778;
   reg _400779_400779 ; 
   reg __400779_400779;
   reg _400780_400780 ; 
   reg __400780_400780;
   reg _400781_400781 ; 
   reg __400781_400781;
   reg _400782_400782 ; 
   reg __400782_400782;
   reg _400783_400783 ; 
   reg __400783_400783;
   reg _400784_400784 ; 
   reg __400784_400784;
   reg _400785_400785 ; 
   reg __400785_400785;
   reg _400786_400786 ; 
   reg __400786_400786;
   reg _400787_400787 ; 
   reg __400787_400787;
   reg _400788_400788 ; 
   reg __400788_400788;
   reg _400789_400789 ; 
   reg __400789_400789;
   reg _400790_400790 ; 
   reg __400790_400790;
   reg _400791_400791 ; 
   reg __400791_400791;
   reg _400792_400792 ; 
   reg __400792_400792;
   reg _400793_400793 ; 
   reg __400793_400793;
   reg _400794_400794 ; 
   reg __400794_400794;
   reg _400795_400795 ; 
   reg __400795_400795;
   reg _400796_400796 ; 
   reg __400796_400796;
   reg _400797_400797 ; 
   reg __400797_400797;
   reg _400798_400798 ; 
   reg __400798_400798;
   reg _400799_400799 ; 
   reg __400799_400799;
   reg _400800_400800 ; 
   reg __400800_400800;
   reg _400801_400801 ; 
   reg __400801_400801;
   reg _400802_400802 ; 
   reg __400802_400802;
   reg _400803_400803 ; 
   reg __400803_400803;
   reg _400804_400804 ; 
   reg __400804_400804;
   reg _400805_400805 ; 
   reg __400805_400805;
   reg _400806_400806 ; 
   reg __400806_400806;
   reg _400807_400807 ; 
   reg __400807_400807;
   reg _400808_400808 ; 
   reg __400808_400808;
   reg _400809_400809 ; 
   reg __400809_400809;
   reg _400810_400810 ; 
   reg __400810_400810;
   reg _400811_400811 ; 
   reg __400811_400811;
   reg _400812_400812 ; 
   reg __400812_400812;
   reg _400813_400813 ; 
   reg __400813_400813;
   reg _400814_400814 ; 
   reg __400814_400814;
   reg _400815_400815 ; 
   reg __400815_400815;
   reg _400816_400816 ; 
   reg __400816_400816;
   reg _400817_400817 ; 
   reg __400817_400817;
   reg _400818_400818 ; 
   reg __400818_400818;
   reg _400819_400819 ; 
   reg __400819_400819;
   reg _400820_400820 ; 
   reg __400820_400820;
   reg _400821_400821 ; 
   reg __400821_400821;
   reg _400822_400822 ; 
   reg __400822_400822;
   reg _400823_400823 ; 
   reg __400823_400823;
   reg _400824_400824 ; 
   reg __400824_400824;
   reg _400825_400825 ; 
   reg __400825_400825;
   reg _400826_400826 ; 
   reg __400826_400826;
   reg _400827_400827 ; 
   reg __400827_400827;
   reg _400828_400828 ; 
   reg __400828_400828;
   reg _400829_400829 ; 
   reg __400829_400829;
   reg _400830_400830 ; 
   reg __400830_400830;
   reg _400831_400831 ; 
   reg __400831_400831;
   reg _400832_400832 ; 
   reg __400832_400832;
   reg _400833_400833 ; 
   reg __400833_400833;
   reg _400834_400834 ; 
   reg __400834_400834;
   reg _400835_400835 ; 
   reg __400835_400835;
   reg _400836_400836 ; 
   reg __400836_400836;
   reg _400837_400837 ; 
   reg __400837_400837;
   reg _400838_400838 ; 
   reg __400838_400838;
   reg _400839_400839 ; 
   reg __400839_400839;
   reg _400840_400840 ; 
   reg __400840_400840;
   reg _400841_400841 ; 
   reg __400841_400841;
   reg _400842_400842 ; 
   reg __400842_400842;
   reg _400843_400843 ; 
   reg __400843_400843;
   reg _400844_400844 ; 
   reg __400844_400844;
   reg _400845_400845 ; 
   reg __400845_400845;
   reg _400846_400846 ; 
   reg __400846_400846;
   reg _400847_400847 ; 
   reg __400847_400847;
   reg _400848_400848 ; 
   reg __400848_400848;
   reg _400849_400849 ; 
   reg __400849_400849;
   reg _400850_400850 ; 
   reg __400850_400850;
   reg _400851_400851 ; 
   reg __400851_400851;
   reg _400852_400852 ; 
   reg __400852_400852;
   reg _400853_400853 ; 
   reg __400853_400853;
   reg _400854_400854 ; 
   reg __400854_400854;
   reg _400855_400855 ; 
   reg __400855_400855;
   reg _400856_400856 ; 
   reg __400856_400856;
   reg _400857_400857 ; 
   reg __400857_400857;
   reg _400858_400858 ; 
   reg __400858_400858;
   reg _400859_400859 ; 
   reg __400859_400859;
   reg _400860_400860 ; 
   reg __400860_400860;
   reg _400861_400861 ; 
   reg __400861_400861;
   reg _400862_400862 ; 
   reg __400862_400862;
   reg _400863_400863 ; 
   reg __400863_400863;
   reg _400864_400864 ; 
   reg __400864_400864;
   reg _400865_400865 ; 
   reg __400865_400865;
   reg _400866_400866 ; 
   reg __400866_400866;
   reg _400867_400867 ; 
   reg __400867_400867;
   reg _400868_400868 ; 
   reg __400868_400868;
   reg _400869_400869 ; 
   reg __400869_400869;
   reg _400870_400870 ; 
   reg __400870_400870;
   reg _400871_400871 ; 
   reg __400871_400871;
   reg _400872_400872 ; 
   reg __400872_400872;
   reg _400873_400873 ; 
   reg __400873_400873;
   reg _400874_400874 ; 
   reg __400874_400874;
   reg _400875_400875 ; 
   reg __400875_400875;
   reg _400876_400876 ; 
   reg __400876_400876;
   reg _400877_400877 ; 
   reg __400877_400877;
   reg _400878_400878 ; 
   reg __400878_400878;
   reg _400879_400879 ; 
   reg __400879_400879;
   reg _400880_400880 ; 
   reg __400880_400880;
   reg _400881_400881 ; 
   reg __400881_400881;
   reg _400882_400882 ; 
   reg __400882_400882;
   reg _400883_400883 ; 
   reg __400883_400883;
   reg _400884_400884 ; 
   reg __400884_400884;
   reg _400885_400885 ; 
   reg __400885_400885;
   reg _400886_400886 ; 
   reg __400886_400886;
   reg _400887_400887 ; 
   reg __400887_400887;
   reg _400888_400888 ; 
   reg __400888_400888;
   reg _400889_400889 ; 
   reg __400889_400889;
   reg _400890_400890 ; 
   reg __400890_400890;
   reg _400891_400891 ; 
   reg __400891_400891;
   reg _400892_400892 ; 
   reg __400892_400892;
   reg _400893_400893 ; 
   reg __400893_400893;
   reg _400894_400894 ; 
   reg __400894_400894;
   reg _400895_400895 ; 
   reg __400895_400895;
   reg _400896_400896 ; 
   reg __400896_400896;
   reg _400897_400897 ; 
   reg __400897_400897;
   reg _400898_400898 ; 
   reg __400898_400898;
   reg _400899_400899 ; 
   reg __400899_400899;
   reg _400900_400900 ; 
   reg __400900_400900;
   reg _400901_400901 ; 
   reg __400901_400901;
   reg _400902_400902 ; 
   reg __400902_400902;
   reg _400903_400903 ; 
   reg __400903_400903;
   reg _400904_400904 ; 
   reg __400904_400904;
   reg _400905_400905 ; 
   reg __400905_400905;
   reg _400906_400906 ; 
   reg __400906_400906;
   reg _400907_400907 ; 
   reg __400907_400907;
   reg _400908_400908 ; 
   reg __400908_400908;
   reg _400909_400909 ; 
   reg __400909_400909;
   reg _400910_400910 ; 
   reg __400910_400910;
   reg _400911_400911 ; 
   reg __400911_400911;
   reg _400912_400912 ; 
   reg __400912_400912;
   reg _400913_400913 ; 
   reg __400913_400913;
   reg _400914_400914 ; 
   reg __400914_400914;
   reg _400915_400915 ; 
   reg __400915_400915;
   reg _400916_400916 ; 
   reg __400916_400916;
   reg _400917_400917 ; 
   reg __400917_400917;
   reg _400918_400918 ; 
   reg __400918_400918;
   reg _400919_400919 ; 
   reg __400919_400919;
   reg _400920_400920 ; 
   reg __400920_400920;
   reg _400921_400921 ; 
   reg __400921_400921;
   reg _400922_400922 ; 
   reg __400922_400922;
   reg _400923_400923 ; 
   reg __400923_400923;
   reg _400924_400924 ; 
   reg __400924_400924;
   reg _400925_400925 ; 
   reg __400925_400925;
   reg _400926_400926 ; 
   reg __400926_400926;
   reg _400927_400927 ; 
   reg __400927_400927;
   reg _400928_400928 ; 
   reg __400928_400928;
   reg _400929_400929 ; 
   reg __400929_400929;
   reg _400930_400930 ; 
   reg __400930_400930;
   reg _400931_400931 ; 
   reg __400931_400931;
   reg _400932_400932 ; 
   reg __400932_400932;
   reg _400933_400933 ; 
   reg __400933_400933;
   reg _400934_400934 ; 
   reg __400934_400934;
   reg _400935_400935 ; 
   reg __400935_400935;
   reg _400936_400936 ; 
   reg __400936_400936;
   reg _400937_400937 ; 
   reg __400937_400937;
   reg _400938_400938 ; 
   reg __400938_400938;
   reg _400939_400939 ; 
   reg __400939_400939;
   reg _400940_400940 ; 
   reg __400940_400940;
   reg _400941_400941 ; 
   reg __400941_400941;
   reg _400942_400942 ; 
   reg __400942_400942;
   reg _400943_400943 ; 
   reg __400943_400943;
   reg _400944_400944 ; 
   reg __400944_400944;
   reg _400945_400945 ; 
   reg __400945_400945;
   reg _400946_400946 ; 
   reg __400946_400946;
   reg _400947_400947 ; 
   reg __400947_400947;
   reg _400948_400948 ; 
   reg __400948_400948;
   reg _400949_400949 ; 
   reg __400949_400949;
   reg _400950_400950 ; 
   reg __400950_400950;
   reg _400951_400951 ; 
   reg __400951_400951;
   reg _400952_400952 ; 
   reg __400952_400952;
   reg _400953_400953 ; 
   reg __400953_400953;
   reg _400954_400954 ; 
   reg __400954_400954;
   reg _400955_400955 ; 
   reg __400955_400955;
   reg _400956_400956 ; 
   reg __400956_400956;
   reg _400957_400957 ; 
   reg __400957_400957;
   reg _400958_400958 ; 
   reg __400958_400958;
   reg _400959_400959 ; 
   reg __400959_400959;
   reg _400960_400960 ; 
   reg __400960_400960;
   reg _400961_400961 ; 
   reg __400961_400961;
   reg _400962_400962 ; 
   reg __400962_400962;
   reg _400963_400963 ; 
   reg __400963_400963;
   reg _400964_400964 ; 
   reg __400964_400964;
   reg _400965_400965 ; 
   reg __400965_400965;
   reg _400966_400966 ; 
   reg __400966_400966;
   reg _400967_400967 ; 
   reg __400967_400967;
   reg _400968_400968 ; 
   reg __400968_400968;
   reg _400969_400969 ; 
   reg __400969_400969;
   reg _400970_400970 ; 
   reg __400970_400970;
   reg _400971_400971 ; 
   reg __400971_400971;
   reg _400972_400972 ; 
   reg __400972_400972;
   reg _400973_400973 ; 
   reg __400973_400973;
   reg _400974_400974 ; 
   reg __400974_400974;
   reg _400975_400975 ; 
   reg __400975_400975;
   reg _400976_400976 ; 
   reg __400976_400976;
   reg _400977_400977 ; 
   reg __400977_400977;
   reg _400978_400978 ; 
   reg __400978_400978;
   reg _400979_400979 ; 
   reg __400979_400979;
   reg _400980_400980 ; 
   reg __400980_400980;
   reg _400981_400981 ; 
   reg __400981_400981;
   reg _400982_400982 ; 
   reg __400982_400982;
   reg _400983_400983 ; 
   reg __400983_400983;
   reg _400984_400984 ; 
   reg __400984_400984;
   reg _400985_400985 ; 
   reg __400985_400985;
   reg _400986_400986 ; 
   reg __400986_400986;
   reg _400987_400987 ; 
   reg __400987_400987;
   reg _400988_400988 ; 
   reg __400988_400988;
   reg _400989_400989 ; 
   reg __400989_400989;
   reg _400990_400990 ; 
   reg __400990_400990;
   reg _400991_400991 ; 
   reg __400991_400991;
   reg _400992_400992 ; 
   reg __400992_400992;
   reg _400993_400993 ; 
   reg __400993_400993;
   reg _400994_400994 ; 
   reg __400994_400994;
   reg _400995_400995 ; 
   reg __400995_400995;
   reg _400996_400996 ; 
   reg __400996_400996;
   reg _400997_400997 ; 
   reg __400997_400997;
   reg _400998_400998 ; 
   reg __400998_400998;
   reg _400999_400999 ; 
   reg __400999_400999;
   reg _401000_401000 ; 
   reg __401000_401000;
   reg _401001_401001 ; 
   reg __401001_401001;
   reg _401002_401002 ; 
   reg __401002_401002;
   reg _401003_401003 ; 
   reg __401003_401003;
   reg _401004_401004 ; 
   reg __401004_401004;
   reg _401005_401005 ; 
   reg __401005_401005;
   reg _401006_401006 ; 
   reg __401006_401006;
   reg _401007_401007 ; 
   reg __401007_401007;
   reg _401008_401008 ; 
   reg __401008_401008;
   reg _401009_401009 ; 
   reg __401009_401009;
   reg _401010_401010 ; 
   reg __401010_401010;
   reg _401011_401011 ; 
   reg __401011_401011;
   reg _401012_401012 ; 
   reg __401012_401012;
   reg _401013_401013 ; 
   reg __401013_401013;
   reg _401014_401014 ; 
   reg __401014_401014;
   reg _401015_401015 ; 
   reg __401015_401015;
   reg _401016_401016 ; 
   reg __401016_401016;
   reg _401017_401017 ; 
   reg __401017_401017;
   reg _401018_401018 ; 
   reg __401018_401018;
   reg _401019_401019 ; 
   reg __401019_401019;
   reg _401020_401020 ; 
   reg __401020_401020;
   reg _401021_401021 ; 
   reg __401021_401021;
   reg _401022_401022 ; 
   reg __401022_401022;
   reg _401023_401023 ; 
   reg __401023_401023;
   reg _401024_401024 ; 
   reg __401024_401024;
   reg _401025_401025 ; 
   reg __401025_401025;
   reg _401026_401026 ; 
   reg __401026_401026;
   reg _401027_401027 ; 
   reg __401027_401027;
   reg _401028_401028 ; 
   reg __401028_401028;
   reg _401029_401029 ; 
   reg __401029_401029;
   reg _401030_401030 ; 
   reg __401030_401030;
   reg _401031_401031 ; 
   reg __401031_401031;
   reg _401032_401032 ; 
   reg __401032_401032;
   reg _401033_401033 ; 
   reg __401033_401033;
   reg _401034_401034 ; 
   reg __401034_401034;
   reg _401035_401035 ; 
   reg __401035_401035;
   reg _401036_401036 ; 
   reg __401036_401036;
   reg _401037_401037 ; 
   reg __401037_401037;
   reg _401038_401038 ; 
   reg __401038_401038;
   reg _401039_401039 ; 
   reg __401039_401039;
   reg _401040_401040 ; 
   reg __401040_401040;
   reg _401041_401041 ; 
   reg __401041_401041;
   reg _401042_401042 ; 
   reg __401042_401042;
   reg _401043_401043 ; 
   reg __401043_401043;
   reg _401044_401044 ; 
   reg __401044_401044;
   reg _401045_401045 ; 
   reg __401045_401045;
   reg _401046_401046 ; 
   reg __401046_401046;
   reg _401047_401047 ; 
   reg __401047_401047;
   reg _401048_401048 ; 
   reg __401048_401048;
   reg _401049_401049 ; 
   reg __401049_401049;
   reg _401050_401050 ; 
   reg __401050_401050;
   reg _401051_401051 ; 
   reg __401051_401051;
   reg _401052_401052 ; 
   reg __401052_401052;
   reg _401053_401053 ; 
   reg __401053_401053;
   reg _401054_401054 ; 
   reg __401054_401054;
   reg _401055_401055 ; 
   reg __401055_401055;
   reg _401056_401056 ; 
   reg __401056_401056;
   reg _401057_401057 ; 
   reg __401057_401057;
   reg _401058_401058 ; 
   reg __401058_401058;
   reg _401059_401059 ; 
   reg __401059_401059;
   reg _401060_401060 ; 
   reg __401060_401060;
   reg _401061_401061 ; 
   reg __401061_401061;
   reg _401062_401062 ; 
   reg __401062_401062;
   reg _401063_401063 ; 
   reg __401063_401063;
   reg _401064_401064 ; 
   reg __401064_401064;
   reg _401065_401065 ; 
   reg __401065_401065;
   reg _401066_401066 ; 
   reg __401066_401066;
   reg _401067_401067 ; 
   reg __401067_401067;
   reg _401068_401068 ; 
   reg __401068_401068;
   reg _401069_401069 ; 
   reg __401069_401069;
   reg _401070_401070 ; 
   reg __401070_401070;
   reg _401071_401071 ; 
   reg __401071_401071;
   reg _401072_401072 ; 
   reg __401072_401072;
   reg _401073_401073 ; 
   reg __401073_401073;
   reg _401074_401074 ; 
   reg __401074_401074;
   reg _401075_401075 ; 
   reg __401075_401075;
   reg _401076_401076 ; 
   reg __401076_401076;
   reg _401077_401077 ; 
   reg __401077_401077;
   reg _401078_401078 ; 
   reg __401078_401078;
   reg _401079_401079 ; 
   reg __401079_401079;
   reg _401080_401080 ; 
   reg __401080_401080;
   reg _401081_401081 ; 
   reg __401081_401081;
   reg _401082_401082 ; 
   reg __401082_401082;
   reg _401083_401083 ; 
   reg __401083_401083;
   reg _401084_401084 ; 
   reg __401084_401084;
   reg _401085_401085 ; 
   reg __401085_401085;
   reg _401086_401086 ; 
   reg __401086_401086;
   reg _401087_401087 ; 
   reg __401087_401087;
   reg _401088_401088 ; 
   reg __401088_401088;
   reg _401089_401089 ; 
   reg __401089_401089;
   reg _401090_401090 ; 
   reg __401090_401090;
   reg _401091_401091 ; 
   reg __401091_401091;
   reg _401092_401092 ; 
   reg __401092_401092;
   reg _401093_401093 ; 
   reg __401093_401093;
   reg _401094_401094 ; 
   reg __401094_401094;
   reg _401095_401095 ; 
   reg __401095_401095;
   reg _401096_401096 ; 
   reg __401096_401096;
   reg _401097_401097 ; 
   reg __401097_401097;
   reg _401098_401098 ; 
   reg __401098_401098;
   reg _401099_401099 ; 
   reg __401099_401099;
   reg _401100_401100 ; 
   reg __401100_401100;
   reg _401101_401101 ; 
   reg __401101_401101;
   reg _401102_401102 ; 
   reg __401102_401102;
   reg _401103_401103 ; 
   reg __401103_401103;
   reg _401104_401104 ; 
   reg __401104_401104;
   reg _401105_401105 ; 
   reg __401105_401105;
   reg _401106_401106 ; 
   reg __401106_401106;
   reg _401107_401107 ; 
   reg __401107_401107;
   reg _401108_401108 ; 
   reg __401108_401108;
   reg _401109_401109 ; 
   reg __401109_401109;
   reg _401110_401110 ; 
   reg __401110_401110;
   reg _401111_401111 ; 
   reg __401111_401111;
   reg _401112_401112 ; 
   reg __401112_401112;
   reg _401113_401113 ; 
   reg __401113_401113;
   reg _401114_401114 ; 
   reg __401114_401114;
   reg _401115_401115 ; 
   reg __401115_401115;
   reg _401116_401116 ; 
   reg __401116_401116;
   reg _401117_401117 ; 
   reg __401117_401117;
   reg _401118_401118 ; 
   reg __401118_401118;
   reg _401119_401119 ; 
   reg __401119_401119;
   reg _401120_401120 ; 
   reg __401120_401120;
   reg _401121_401121 ; 
   reg __401121_401121;
   reg _401122_401122 ; 
   reg __401122_401122;
   reg _401123_401123 ; 
   reg __401123_401123;
   reg _401124_401124 ; 
   reg __401124_401124;
   reg _401125_401125 ; 
   reg __401125_401125;
   reg _401126_401126 ; 
   reg __401126_401126;
   reg _401127_401127 ; 
   reg __401127_401127;
   reg _401128_401128 ; 
   reg __401128_401128;
   reg _401129_401129 ; 
   reg __401129_401129;
   reg _401130_401130 ; 
   reg __401130_401130;
   reg _401131_401131 ; 
   reg __401131_401131;
   reg _401132_401132 ; 
   reg __401132_401132;
   reg _401133_401133 ; 
   reg __401133_401133;
   reg _401134_401134 ; 
   reg __401134_401134;
   reg _401135_401135 ; 
   reg __401135_401135;
   reg _401136_401136 ; 
   reg __401136_401136;
   reg _401137_401137 ; 
   reg __401137_401137;
   reg _401138_401138 ; 
   reg __401138_401138;
   reg _401139_401139 ; 
   reg __401139_401139;
   reg _401140_401140 ; 
   reg __401140_401140;
   reg _401141_401141 ; 
   reg __401141_401141;
   reg _401142_401142 ; 
   reg __401142_401142;
   reg _401143_401143 ; 
   reg __401143_401143;
   reg _401144_401144 ; 
   reg __401144_401144;
   reg _401145_401145 ; 
   reg __401145_401145;
   reg _401146_401146 ; 
   reg __401146_401146;
   reg _401147_401147 ; 
   reg __401147_401147;
   reg _401148_401148 ; 
   reg __401148_401148;
   reg _401149_401149 ; 
   reg __401149_401149;
   reg _401150_401150 ; 
   reg __401150_401150;
   reg _401151_401151 ; 
   reg __401151_401151;
   reg _401152_401152 ; 
   reg __401152_401152;
   reg _401153_401153 ; 
   reg __401153_401153;
   reg _401154_401154 ; 
   reg __401154_401154;
   reg _401155_401155 ; 
   reg __401155_401155;
   reg _401156_401156 ; 
   reg __401156_401156;
   reg _401157_401157 ; 
   reg __401157_401157;
   reg _401158_401158 ; 
   reg __401158_401158;
   reg _401159_401159 ; 
   reg __401159_401159;
   reg _401160_401160 ; 
   reg __401160_401160;
   reg _401161_401161 ; 
   reg __401161_401161;
   reg _401162_401162 ; 
   reg __401162_401162;
   reg _401163_401163 ; 
   reg __401163_401163;
   reg _401164_401164 ; 
   reg __401164_401164;
   reg _401165_401165 ; 
   reg __401165_401165;
   reg _401166_401166 ; 
   reg __401166_401166;
   reg _401167_401167 ; 
   reg __401167_401167;
   reg _401168_401168 ; 
   reg __401168_401168;
   reg _401169_401169 ; 
   reg __401169_401169;
   reg _401170_401170 ; 
   reg __401170_401170;
   reg _401171_401171 ; 
   reg __401171_401171;
   reg _401172_401172 ; 
   reg __401172_401172;
   reg _401173_401173 ; 
   reg __401173_401173;
   reg _401174_401174 ; 
   reg __401174_401174;
   reg _401175_401175 ; 
   reg __401175_401175;
   reg _401176_401176 ; 
   reg __401176_401176;
   reg _401177_401177 ; 
   reg __401177_401177;
   reg _401178_401178 ; 
   reg __401178_401178;
   reg _401179_401179 ; 
   reg __401179_401179;
   reg _401180_401180 ; 
   reg __401180_401180;
   reg _401181_401181 ; 
   reg __401181_401181;
   reg _401182_401182 ; 
   reg __401182_401182;
   reg _401183_401183 ; 
   reg __401183_401183;
   reg _401184_401184 ; 
   reg __401184_401184;
   reg _401185_401185 ; 
   reg __401185_401185;
   reg _401186_401186 ; 
   reg __401186_401186;
   reg _401187_401187 ; 
   reg __401187_401187;
   reg _401188_401188 ; 
   reg __401188_401188;
   reg _401189_401189 ; 
   reg __401189_401189;
   reg _401190_401190 ; 
   reg __401190_401190;
   reg _401191_401191 ; 
   reg __401191_401191;
   reg _401192_401192 ; 
   reg __401192_401192;
   reg _401193_401193 ; 
   reg __401193_401193;
   reg _401194_401194 ; 
   reg __401194_401194;
   reg _401195_401195 ; 
   reg __401195_401195;
   reg _401196_401196 ; 
   reg __401196_401196;
   reg _401197_401197 ; 
   reg __401197_401197;
   reg _401198_401198 ; 
   reg __401198_401198;
   reg _401199_401199 ; 
   reg __401199_401199;
   reg _401200_401200 ; 
   reg __401200_401200;
   reg _401201_401201 ; 
   reg __401201_401201;
   reg _401202_401202 ; 
   reg __401202_401202;
   reg _401203_401203 ; 
   reg __401203_401203;
   reg _401204_401204 ; 
   reg __401204_401204;
   reg _401205_401205 ; 
   reg __401205_401205;
   reg _401206_401206 ; 
   reg __401206_401206;
   reg _401207_401207 ; 
   reg __401207_401207;
   reg _401208_401208 ; 
   reg __401208_401208;
   reg _401209_401209 ; 
   reg __401209_401209;
   reg _401210_401210 ; 
   reg __401210_401210;
   reg _401211_401211 ; 
   reg __401211_401211;
   reg _401212_401212 ; 
   reg __401212_401212;
   reg _401213_401213 ; 
   reg __401213_401213;
   reg _401214_401214 ; 
   reg __401214_401214;
   reg _401215_401215 ; 
   reg __401215_401215;
   reg _401216_401216 ; 
   reg __401216_401216;
   reg _401217_401217 ; 
   reg __401217_401217;
   reg _401218_401218 ; 
   reg __401218_401218;
   reg _401219_401219 ; 
   reg __401219_401219;
   reg _401220_401220 ; 
   reg __401220_401220;
   reg _401221_401221 ; 
   reg __401221_401221;
   reg _401222_401222 ; 
   reg __401222_401222;
   reg _401223_401223 ; 
   reg __401223_401223;
   reg _401224_401224 ; 
   reg __401224_401224;
   reg _401225_401225 ; 
   reg __401225_401225;
   reg _401226_401226 ; 
   reg __401226_401226;
   reg _401227_401227 ; 
   reg __401227_401227;
   reg _401228_401228 ; 
   reg __401228_401228;
   reg _401229_401229 ; 
   reg __401229_401229;
   reg _401230_401230 ; 
   reg __401230_401230;
   reg _401231_401231 ; 
   reg __401231_401231;
   reg _401232_401232 ; 
   reg __401232_401232;
   reg _401233_401233 ; 
   reg __401233_401233;
   reg _401234_401234 ; 
   reg __401234_401234;
   reg _401235_401235 ; 
   reg __401235_401235;
   reg _401236_401236 ; 
   reg __401236_401236;
   reg _401237_401237 ; 
   reg __401237_401237;
   reg _401238_401238 ; 
   reg __401238_401238;
   reg _401239_401239 ; 
   reg __401239_401239;
   reg _401240_401240 ; 
   reg __401240_401240;
   reg _401241_401241 ; 
   reg __401241_401241;
   reg _401242_401242 ; 
   reg __401242_401242;
   reg _401243_401243 ; 
   reg __401243_401243;
   reg _401244_401244 ; 
   reg __401244_401244;
   reg _401245_401245 ; 
   reg __401245_401245;
   reg _401246_401246 ; 
   reg __401246_401246;
   reg _401247_401247 ; 
   reg __401247_401247;
   reg _401248_401248 ; 
   reg __401248_401248;
   reg _401249_401249 ; 
   reg __401249_401249;
   reg _401250_401250 ; 
   reg __401250_401250;
   reg _401251_401251 ; 
   reg __401251_401251;
   reg _401252_401252 ; 
   reg __401252_401252;
   reg _401253_401253 ; 
   reg __401253_401253;
   reg _401254_401254 ; 
   reg __401254_401254;
   reg _401255_401255 ; 
   reg __401255_401255;
   reg _401256_401256 ; 
   reg __401256_401256;
   reg _401257_401257 ; 
   reg __401257_401257;
   reg _401258_401258 ; 
   reg __401258_401258;
   reg _401259_401259 ; 
   reg __401259_401259;
   reg _401260_401260 ; 
   reg __401260_401260;
   reg _401261_401261 ; 
   reg __401261_401261;
   reg _401262_401262 ; 
   reg __401262_401262;
   reg _401263_401263 ; 
   reg __401263_401263;
   reg _401264_401264 ; 
   reg __401264_401264;
   reg _401265_401265 ; 
   reg __401265_401265;
   reg _401266_401266 ; 
   reg __401266_401266;
   reg _401267_401267 ; 
   reg __401267_401267;
   reg _401268_401268 ; 
   reg __401268_401268;
   reg _401269_401269 ; 
   reg __401269_401269;
   reg _401270_401270 ; 
   reg __401270_401270;
   reg _401271_401271 ; 
   reg __401271_401271;
   reg _401272_401272 ; 
   reg __401272_401272;
   reg _401273_401273 ; 
   reg __401273_401273;
   reg _401274_401274 ; 
   reg __401274_401274;
   reg _401275_401275 ; 
   reg __401275_401275;
   reg _401276_401276 ; 
   reg __401276_401276;
   reg _401277_401277 ; 
   reg __401277_401277;
   reg _401278_401278 ; 
   reg __401278_401278;
   reg _401279_401279 ; 
   reg __401279_401279;
   reg _401280_401280 ; 
   reg __401280_401280;
   reg _401281_401281 ; 
   reg __401281_401281;
   reg _401282_401282 ; 
   reg __401282_401282;
   reg _401283_401283 ; 
   reg __401283_401283;
   reg _401284_401284 ; 
   reg __401284_401284;
   reg _401285_401285 ; 
   reg __401285_401285;
   reg _401286_401286 ; 
   reg __401286_401286;
   reg _401287_401287 ; 
   reg __401287_401287;
   reg _401288_401288 ; 
   reg __401288_401288;
   reg _401289_401289 ; 
   reg __401289_401289;
   reg _401290_401290 ; 
   reg __401290_401290;
   reg _401291_401291 ; 
   reg __401291_401291;
   reg _401292_401292 ; 
   reg __401292_401292;
   reg _401293_401293 ; 
   reg __401293_401293;
   reg _401294_401294 ; 
   reg __401294_401294;
   reg _401295_401295 ; 
   reg __401295_401295;
   reg _401296_401296 ; 
   reg __401296_401296;
   reg _401297_401297 ; 
   reg __401297_401297;
   reg _401298_401298 ; 
   reg __401298_401298;
   reg _401299_401299 ; 
   reg __401299_401299;
   reg _401300_401300 ; 
   reg __401300_401300;
   reg _401301_401301 ; 
   reg __401301_401301;
   reg _401302_401302 ; 
   reg __401302_401302;
   reg _401303_401303 ; 
   reg __401303_401303;
   reg _401304_401304 ; 
   reg __401304_401304;
   reg _401305_401305 ; 
   reg __401305_401305;
   reg _401306_401306 ; 
   reg __401306_401306;
   reg _401307_401307 ; 
   reg __401307_401307;
   reg _401308_401308 ; 
   reg __401308_401308;
   reg _401309_401309 ; 
   reg __401309_401309;
   reg _401310_401310 ; 
   reg __401310_401310;
   reg _401311_401311 ; 
   reg __401311_401311;
   reg _401312_401312 ; 
   reg __401312_401312;
   reg _401313_401313 ; 
   reg __401313_401313;
   reg _401314_401314 ; 
   reg __401314_401314;
   reg _401315_401315 ; 
   reg __401315_401315;
   reg _401316_401316 ; 
   reg __401316_401316;
   reg _401317_401317 ; 
   reg __401317_401317;
   reg _401318_401318 ; 
   reg __401318_401318;
   reg _401319_401319 ; 
   reg __401319_401319;
   reg _401320_401320 ; 
   reg __401320_401320;
   reg _401321_401321 ; 
   reg __401321_401321;
   reg _401322_401322 ; 
   reg __401322_401322;
   reg _401323_401323 ; 
   reg __401323_401323;
   reg _401324_401324 ; 
   reg __401324_401324;
   reg _401325_401325 ; 
   reg __401325_401325;
   reg _401326_401326 ; 
   reg __401326_401326;
   reg _401327_401327 ; 
   reg __401327_401327;
   reg _401328_401328 ; 
   reg __401328_401328;
   reg _401329_401329 ; 
   reg __401329_401329;
   reg _401330_401330 ; 
   reg __401330_401330;
   reg _401331_401331 ; 
   reg __401331_401331;
   reg _401332_401332 ; 
   reg __401332_401332;
   reg _401333_401333 ; 
   reg __401333_401333;
   reg _401334_401334 ; 
   reg __401334_401334;
   reg _401335_401335 ; 
   reg __401335_401335;
   reg _401336_401336 ; 
   reg __401336_401336;
   reg _401337_401337 ; 
   reg __401337_401337;
   reg _401338_401338 ; 
   reg __401338_401338;
   reg _401339_401339 ; 
   reg __401339_401339;
   reg _401340_401340 ; 
   reg __401340_401340;
   reg _401341_401341 ; 
   reg __401341_401341;
   reg _401342_401342 ; 
   reg __401342_401342;
   reg _401343_401343 ; 
   reg __401343_401343;
   reg _401344_401344 ; 
   reg __401344_401344;
   reg _401345_401345 ; 
   reg __401345_401345;
   reg _401346_401346 ; 
   reg __401346_401346;
   reg _401347_401347 ; 
   reg __401347_401347;
   reg _401348_401348 ; 
   reg __401348_401348;
   reg _401349_401349 ; 
   reg __401349_401349;
   reg _401350_401350 ; 
   reg __401350_401350;
   reg _401351_401351 ; 
   reg __401351_401351;
   reg _401352_401352 ; 
   reg __401352_401352;
   reg _401353_401353 ; 
   reg __401353_401353;
   reg _401354_401354 ; 
   reg __401354_401354;
   reg _401355_401355 ; 
   reg __401355_401355;
   reg _401356_401356 ; 
   reg __401356_401356;
   reg _401357_401357 ; 
   reg __401357_401357;
   reg _401358_401358 ; 
   reg __401358_401358;
   reg _401359_401359 ; 
   reg __401359_401359;
   reg _401360_401360 ; 
   reg __401360_401360;
   reg _401361_401361 ; 
   reg __401361_401361;
   reg _401362_401362 ; 
   reg __401362_401362;
   reg _401363_401363 ; 
   reg __401363_401363;
   reg _401364_401364 ; 
   reg __401364_401364;
   reg _401365_401365 ; 
   reg __401365_401365;
   reg _401366_401366 ; 
   reg __401366_401366;
   reg _401367_401367 ; 
   reg __401367_401367;
   reg _401368_401368 ; 
   reg __401368_401368;
   reg _401369_401369 ; 
   reg __401369_401369;
   reg _401370_401370 ; 
   reg __401370_401370;
   reg _401371_401371 ; 
   reg __401371_401371;
   reg _401372_401372 ; 
   reg __401372_401372;
   reg _401373_401373 ; 
   reg __401373_401373;
   reg _401374_401374 ; 
   reg __401374_401374;
   reg _401375_401375 ; 
   reg __401375_401375;
   reg _401376_401376 ; 
   reg __401376_401376;
   reg _401377_401377 ; 
   reg __401377_401377;
   reg _401378_401378 ; 
   reg __401378_401378;
   reg _401379_401379 ; 
   reg __401379_401379;
   reg _401380_401380 ; 
   reg __401380_401380;
   reg _401381_401381 ; 
   reg __401381_401381;
   reg _401382_401382 ; 
   reg __401382_401382;
   reg _401383_401383 ; 
   reg __401383_401383;
   reg _401384_401384 ; 
   reg __401384_401384;
   reg _401385_401385 ; 
   reg __401385_401385;
   reg _401386_401386 ; 
   reg __401386_401386;
   reg _401387_401387 ; 
   reg __401387_401387;
   reg _401388_401388 ; 
   reg __401388_401388;
   reg _401389_401389 ; 
   reg __401389_401389;
   reg _401390_401390 ; 
   reg __401390_401390;
   reg _401391_401391 ; 
   reg __401391_401391;
   reg _401392_401392 ; 
   reg __401392_401392;
   reg _401393_401393 ; 
   reg __401393_401393;
   reg _401394_401394 ; 
   reg __401394_401394;
   reg _401395_401395 ; 
   reg __401395_401395;
   reg _401396_401396 ; 
   reg __401396_401396;
   reg _401397_401397 ; 
   reg __401397_401397;
   reg _401398_401398 ; 
   reg __401398_401398;
   reg _401399_401399 ; 
   reg __401399_401399;
   reg _401400_401400 ; 
   reg __401400_401400;
   reg _401401_401401 ; 
   reg __401401_401401;
   reg _401402_401402 ; 
   reg __401402_401402;
   reg _401403_401403 ; 
   reg __401403_401403;
   reg _401404_401404 ; 
   reg __401404_401404;
   reg _401405_401405 ; 
   reg __401405_401405;
   reg _401406_401406 ; 
   reg __401406_401406;
   reg _401407_401407 ; 
   reg __401407_401407;
   reg _401408_401408 ; 
   reg __401408_401408;
   reg _401409_401409 ; 
   reg __401409_401409;
   reg _401410_401410 ; 
   reg __401410_401410;
   reg _401411_401411 ; 
   reg __401411_401411;
   reg _401412_401412 ; 
   reg __401412_401412;
   reg _401413_401413 ; 
   reg __401413_401413;
   reg _401414_401414 ; 
   reg __401414_401414;
   reg _401415_401415 ; 
   reg __401415_401415;
   reg _401416_401416 ; 
   reg __401416_401416;
   reg _401417_401417 ; 
   reg __401417_401417;
   reg _401418_401418 ; 
   reg __401418_401418;
   reg _401419_401419 ; 
   reg __401419_401419;
   reg _401420_401420 ; 
   reg __401420_401420;
   reg _401421_401421 ; 
   reg __401421_401421;
   reg _401422_401422 ; 
   reg __401422_401422;
   reg _401423_401423 ; 
   reg __401423_401423;
   reg _401424_401424 ; 
   reg __401424_401424;
   reg _401425_401425 ; 
   reg __401425_401425;
   reg _401426_401426 ; 
   reg __401426_401426;
   reg _401427_401427 ; 
   reg __401427_401427;
   reg _401428_401428 ; 
   reg __401428_401428;
   reg _401429_401429 ; 
   reg __401429_401429;
   reg _401430_401430 ; 
   reg __401430_401430;
   reg _401431_401431 ; 
   reg __401431_401431;
   reg _401432_401432 ; 
   reg __401432_401432;
   reg _401433_401433 ; 
   reg __401433_401433;
   reg _401434_401434 ; 
   reg __401434_401434;
   reg _401435_401435 ; 
   reg __401435_401435;
   reg _401436_401436 ; 
   reg __401436_401436;
   reg _401437_401437 ; 
   reg __401437_401437;
   reg _401438_401438 ; 
   reg __401438_401438;
   reg _401439_401439 ; 
   reg __401439_401439;
   reg _401440_401440 ; 
   reg __401440_401440;
   reg _401441_401441 ; 
   reg __401441_401441;
   reg _401442_401442 ; 
   reg __401442_401442;
   reg _401443_401443 ; 
   reg __401443_401443;
   reg _401444_401444 ; 
   reg __401444_401444;
   reg _401445_401445 ; 
   reg __401445_401445;
   reg _401446_401446 ; 
   reg __401446_401446;
   reg _401447_401447 ; 
   reg __401447_401447;
   reg _401448_401448 ; 
   reg __401448_401448;
   reg _401449_401449 ; 
   reg __401449_401449;
   reg _401450_401450 ; 
   reg __401450_401450;
   reg _401451_401451 ; 
   reg __401451_401451;
   reg _401452_401452 ; 
   reg __401452_401452;
   reg _401453_401453 ; 
   reg __401453_401453;
   reg _401454_401454 ; 
   reg __401454_401454;
   reg _401455_401455 ; 
   reg __401455_401455;
   reg _401456_401456 ; 
   reg __401456_401456;
   reg _401457_401457 ; 
   reg __401457_401457;
   reg _401458_401458 ; 
   reg __401458_401458;
   reg _401459_401459 ; 
   reg __401459_401459;
   reg _401460_401460 ; 
   reg __401460_401460;
   reg _401461_401461 ; 
   reg __401461_401461;
   reg _401462_401462 ; 
   reg __401462_401462;
   reg _401463_401463 ; 
   reg __401463_401463;
   reg _401464_401464 ; 
   reg __401464_401464;
   reg _401465_401465 ; 
   reg __401465_401465;
   reg _401466_401466 ; 
   reg __401466_401466;
   reg _401467_401467 ; 
   reg __401467_401467;
   reg _401468_401468 ; 
   reg __401468_401468;
   reg _401469_401469 ; 
   reg __401469_401469;
   reg _401470_401470 ; 
   reg __401470_401470;
   reg _401471_401471 ; 
   reg __401471_401471;
   reg _401472_401472 ; 
   reg __401472_401472;
   reg _401473_401473 ; 
   reg __401473_401473;
   reg _401474_401474 ; 
   reg __401474_401474;
   reg _401475_401475 ; 
   reg __401475_401475;
   reg _401476_401476 ; 
   reg __401476_401476;
   reg _401477_401477 ; 
   reg __401477_401477;
   reg _401478_401478 ; 
   reg __401478_401478;
   reg _401479_401479 ; 
   reg __401479_401479;
   reg _401480_401480 ; 
   reg __401480_401480;
   reg _401481_401481 ; 
   reg __401481_401481;
   reg _401482_401482 ; 
   reg __401482_401482;
   reg _401483_401483 ; 
   reg __401483_401483;
   reg _401484_401484 ; 
   reg __401484_401484;
   reg _401485_401485 ; 
   reg __401485_401485;
   reg _401486_401486 ; 
   reg __401486_401486;
   reg _401487_401487 ; 
   reg __401487_401487;
   reg _401488_401488 ; 
   reg __401488_401488;
   reg _401489_401489 ; 
   reg __401489_401489;
   reg _401490_401490 ; 
   reg __401490_401490;
   reg _401491_401491 ; 
   reg __401491_401491;
   reg _401492_401492 ; 
   reg __401492_401492;
   reg _401493_401493 ; 
   reg __401493_401493;
   reg _401494_401494 ; 
   reg __401494_401494;
   reg _401495_401495 ; 
   reg __401495_401495;
   reg _401496_401496 ; 
   reg __401496_401496;
   reg _401497_401497 ; 
   reg __401497_401497;
   reg _401498_401498 ; 
   reg __401498_401498;
   reg _401499_401499 ; 
   reg __401499_401499;
   reg _401500_401500 ; 
   reg __401500_401500;
   reg _401501_401501 ; 
   reg __401501_401501;
   reg _401502_401502 ; 
   reg __401502_401502;
   reg _401503_401503 ; 
   reg __401503_401503;
   reg _401504_401504 ; 
   reg __401504_401504;
   reg _401505_401505 ; 
   reg __401505_401505;
   reg _401506_401506 ; 
   reg __401506_401506;
   reg _401507_401507 ; 
   reg __401507_401507;
   reg _401508_401508 ; 
   reg __401508_401508;
   reg _401509_401509 ; 
   reg __401509_401509;
   reg _401510_401510 ; 
   reg __401510_401510;
   reg _401511_401511 ; 
   reg __401511_401511;
   reg _401512_401512 ; 
   reg __401512_401512;
   reg _401513_401513 ; 
   reg __401513_401513;
   reg _401514_401514 ; 
   reg __401514_401514;
   reg _401515_401515 ; 
   reg __401515_401515;
   reg _401516_401516 ; 
   reg __401516_401516;
   reg _401517_401517 ; 
   reg __401517_401517;
   reg _401518_401518 ; 
   reg __401518_401518;
   reg _401519_401519 ; 
   reg __401519_401519;
   reg _401520_401520 ; 
   reg __401520_401520;
   reg _401521_401521 ; 
   reg __401521_401521;
   reg _401522_401522 ; 
   reg __401522_401522;
   reg _401523_401523 ; 
   reg __401523_401523;
   reg _401524_401524 ; 
   reg __401524_401524;
   reg _401525_401525 ; 
   reg __401525_401525;
   reg _401526_401526 ; 
   reg __401526_401526;
   reg _401527_401527 ; 
   reg __401527_401527;
   reg _401528_401528 ; 
   reg __401528_401528;
   reg _401529_401529 ; 
   reg __401529_401529;
   reg _401530_401530 ; 
   reg __401530_401530;
   reg _401531_401531 ; 
   reg __401531_401531;
   reg _401532_401532 ; 
   reg __401532_401532;
   reg _401533_401533 ; 
   reg __401533_401533;
   reg _401534_401534 ; 
   reg __401534_401534;
   reg _401535_401535 ; 
   reg __401535_401535;
   reg _401536_401536 ; 
   reg __401536_401536;
   reg _401537_401537 ; 
   reg __401537_401537;
   reg _401538_401538 ; 
   reg __401538_401538;
   reg _401539_401539 ; 
   reg __401539_401539;
   reg _401540_401540 ; 
   reg __401540_401540;
   reg _401541_401541 ; 
   reg __401541_401541;
   reg _401542_401542 ; 
   reg __401542_401542;
   reg _401543_401543 ; 
   reg __401543_401543;
   reg _401544_401544 ; 
   reg __401544_401544;
   reg _401545_401545 ; 
   reg __401545_401545;
   reg _401546_401546 ; 
   reg __401546_401546;
   reg _401547_401547 ; 
   reg __401547_401547;
   reg _401548_401548 ; 
   reg __401548_401548;
   reg _401549_401549 ; 
   reg __401549_401549;
   reg _401550_401550 ; 
   reg __401550_401550;
   reg _401551_401551 ; 
   reg __401551_401551;
   reg _401552_401552 ; 
   reg __401552_401552;
   reg _401553_401553 ; 
   reg __401553_401553;
   reg _401554_401554 ; 
   reg __401554_401554;
   reg _401555_401555 ; 
   reg __401555_401555;
   reg _401556_401556 ; 
   reg __401556_401556;
   reg _401557_401557 ; 
   reg __401557_401557;
   reg _401558_401558 ; 
   reg __401558_401558;
   reg _401559_401559 ; 
   reg __401559_401559;
   reg _401560_401560 ; 
   reg __401560_401560;
   reg _401561_401561 ; 
   reg __401561_401561;
   reg _401562_401562 ; 
   reg __401562_401562;
   reg _401563_401563 ; 
   reg __401563_401563;
   reg _401564_401564 ; 
   reg __401564_401564;
   reg _401565_401565 ; 
   reg __401565_401565;
   reg _401566_401566 ; 
   reg __401566_401566;
   reg _401567_401567 ; 
   reg __401567_401567;
   reg _401568_401568 ; 
   reg __401568_401568;
   reg _401569_401569 ; 
   reg __401569_401569;
   reg _401570_401570 ; 
   reg __401570_401570;
   reg _401571_401571 ; 
   reg __401571_401571;
   reg _401572_401572 ; 
   reg __401572_401572;
   reg _401573_401573 ; 
   reg __401573_401573;
   reg _401574_401574 ; 
   reg __401574_401574;
   reg _401575_401575 ; 
   reg __401575_401575;
   reg _401576_401576 ; 
   reg __401576_401576;
   reg _401577_401577 ; 
   reg __401577_401577;
   reg _401578_401578 ; 
   reg __401578_401578;
   reg _401579_401579 ; 
   reg __401579_401579;
   reg _401580_401580 ; 
   reg __401580_401580;
   reg _401581_401581 ; 
   reg __401581_401581;
   reg _401582_401582 ; 
   reg __401582_401582;
   reg _401583_401583 ; 
   reg __401583_401583;
   reg _401584_401584 ; 
   reg __401584_401584;
   reg _401585_401585 ; 
   reg __401585_401585;
   reg _401586_401586 ; 
   reg __401586_401586;
   reg _401587_401587 ; 
   reg __401587_401587;
   reg _401588_401588 ; 
   reg __401588_401588;
   reg _401589_401589 ; 
   reg __401589_401589;
   reg _401590_401590 ; 
   reg __401590_401590;
   reg _401591_401591 ; 
   reg __401591_401591;
   reg _401592_401592 ; 
   reg __401592_401592;
   reg _401593_401593 ; 
   reg __401593_401593;
   reg _401594_401594 ; 
   reg __401594_401594;
   reg _401595_401595 ; 
   reg __401595_401595;
   reg _401596_401596 ; 
   reg __401596_401596;
   reg _401597_401597 ; 
   reg __401597_401597;
   reg _401598_401598 ; 
   reg __401598_401598;
   reg _401599_401599 ; 
   reg __401599_401599;
   reg _401600_401600 ; 
   reg __401600_401600;
   reg _401601_401601 ; 
   reg __401601_401601;
   reg _401602_401602 ; 
   reg __401602_401602;
   reg _401603_401603 ; 
   reg __401603_401603;
   reg _401604_401604 ; 
   reg __401604_401604;
   reg _401605_401605 ; 
   reg __401605_401605;
   reg _401606_401606 ; 
   reg __401606_401606;
   reg _401607_401607 ; 
   reg __401607_401607;
   reg _401608_401608 ; 
   reg __401608_401608;
   reg _401609_401609 ; 
   reg __401609_401609;
   reg _401610_401610 ; 
   reg __401610_401610;
   reg _401611_401611 ; 
   reg __401611_401611;
   reg _401612_401612 ; 
   reg __401612_401612;
   reg _401613_401613 ; 
   reg __401613_401613;
   reg _401614_401614 ; 
   reg __401614_401614;
   reg _401615_401615 ; 
   reg __401615_401615;
   reg _401616_401616 ; 
   reg __401616_401616;
   reg _401617_401617 ; 
   reg __401617_401617;
   reg _401618_401618 ; 
   reg __401618_401618;
   reg _401619_401619 ; 
   reg __401619_401619;
   reg _401620_401620 ; 
   reg __401620_401620;
   reg _401621_401621 ; 
   reg __401621_401621;
   reg _401622_401622 ; 
   reg __401622_401622;
   reg _401623_401623 ; 
   reg __401623_401623;
   reg _401624_401624 ; 
   reg __401624_401624;
   reg _401625_401625 ; 
   reg __401625_401625;
   reg _401626_401626 ; 
   reg __401626_401626;
   reg _401627_401627 ; 
   reg __401627_401627;
   reg _401628_401628 ; 
   reg __401628_401628;
   reg _401629_401629 ; 
   reg __401629_401629;
   reg _401630_401630 ; 
   reg __401630_401630;
   reg _401631_401631 ; 
   reg __401631_401631;
   reg _401632_401632 ; 
   reg __401632_401632;
   reg _401633_401633 ; 
   reg __401633_401633;
   reg _401634_401634 ; 
   reg __401634_401634;
   reg _401635_401635 ; 
   reg __401635_401635;
   reg _401636_401636 ; 
   reg __401636_401636;
   reg _401637_401637 ; 
   reg __401637_401637;
   reg _401638_401638 ; 
   reg __401638_401638;
   reg _401639_401639 ; 
   reg __401639_401639;
   reg _401640_401640 ; 
   reg __401640_401640;
   reg _401641_401641 ; 
   reg __401641_401641;
   reg _401642_401642 ; 
   reg __401642_401642;
   reg _401643_401643 ; 
   reg __401643_401643;
   reg _401644_401644 ; 
   reg __401644_401644;
   reg _401645_401645 ; 
   reg __401645_401645;
   reg _401646_401646 ; 
   reg __401646_401646;
   reg _401647_401647 ; 
   reg __401647_401647;
   reg _401648_401648 ; 
   reg __401648_401648;
   reg _401649_401649 ; 
   reg __401649_401649;
   reg _401650_401650 ; 
   reg __401650_401650;
   reg _401651_401651 ; 
   reg __401651_401651;
   reg _401652_401652 ; 
   reg __401652_401652;
   reg _401653_401653 ; 
   reg __401653_401653;
   reg _401654_401654 ; 
   reg __401654_401654;
   reg _401655_401655 ; 
   reg __401655_401655;
   reg _401656_401656 ; 
   reg __401656_401656;
   reg _401657_401657 ; 
   reg __401657_401657;
   reg _401658_401658 ; 
   reg __401658_401658;
   reg _401659_401659 ; 
   reg __401659_401659;
   reg _401660_401660 ; 
   reg __401660_401660;
   reg _401661_401661 ; 
   reg __401661_401661;
   reg _401662_401662 ; 
   reg __401662_401662;
   reg _401663_401663 ; 
   reg __401663_401663;
   reg _401664_401664 ; 
   reg __401664_401664;
   reg _401665_401665 ; 
   reg __401665_401665;
   reg _401666_401666 ; 
   reg __401666_401666;
   reg _401667_401667 ; 
   reg __401667_401667;
   reg _401668_401668 ; 
   reg __401668_401668;
   reg _401669_401669 ; 
   reg __401669_401669;
   reg _401670_401670 ; 
   reg __401670_401670;
   reg _401671_401671 ; 
   reg __401671_401671;
   reg _401672_401672 ; 
   reg __401672_401672;
   reg _401673_401673 ; 
   reg __401673_401673;
   reg _401674_401674 ; 
   reg __401674_401674;
   reg _401675_401675 ; 
   reg __401675_401675;
   reg _401676_401676 ; 
   reg __401676_401676;
   reg _401677_401677 ; 
   reg __401677_401677;
   reg _401678_401678 ; 
   reg __401678_401678;
   reg _401679_401679 ; 
   reg __401679_401679;
   reg _401680_401680 ; 
   reg __401680_401680;
   reg _401681_401681 ; 
   reg __401681_401681;
   reg _401682_401682 ; 
   reg __401682_401682;
   reg _401683_401683 ; 
   reg __401683_401683;
   reg _401684_401684 ; 
   reg __401684_401684;
   reg _401685_401685 ; 
   reg __401685_401685;
   reg _401686_401686 ; 
   reg __401686_401686;
   reg _401687_401687 ; 
   reg __401687_401687;
   reg _401688_401688 ; 
   reg __401688_401688;
   reg _401689_401689 ; 
   reg __401689_401689;
   reg _401690_401690 ; 
   reg __401690_401690;
   reg _401691_401691 ; 
   reg __401691_401691;
   reg _401692_401692 ; 
   reg __401692_401692;
   reg _401693_401693 ; 
   reg __401693_401693;
   reg _401694_401694 ; 
   reg __401694_401694;
   reg _401695_401695 ; 
   reg __401695_401695;
   reg _401696_401696 ; 
   reg __401696_401696;
   reg _401697_401697 ; 
   reg __401697_401697;
   reg _401698_401698 ; 
   reg __401698_401698;
   reg _401699_401699 ; 
   reg __401699_401699;
   reg _401700_401700 ; 
   reg __401700_401700;
   reg _401701_401701 ; 
   reg __401701_401701;
   reg _401702_401702 ; 
   reg __401702_401702;
   reg _401703_401703 ; 
   reg __401703_401703;
   reg _401704_401704 ; 
   reg __401704_401704;
   reg _401705_401705 ; 
   reg __401705_401705;
   reg _401706_401706 ; 
   reg __401706_401706;
   reg _401707_401707 ; 
   reg __401707_401707;
   reg _401708_401708 ; 
   reg __401708_401708;
   reg _401709_401709 ; 
   reg __401709_401709;
   reg _401710_401710 ; 
   reg __401710_401710;
   reg _401711_401711 ; 
   reg __401711_401711;
   reg _401712_401712 ; 
   reg __401712_401712;
   reg _401713_401713 ; 
   reg __401713_401713;
   reg _401714_401714 ; 
   reg __401714_401714;
   reg _401715_401715 ; 
   reg __401715_401715;
   reg _401716_401716 ; 
   reg __401716_401716;
   reg _401717_401717 ; 
   reg __401717_401717;
   reg _401718_401718 ; 
   reg __401718_401718;
   reg _401719_401719 ; 
   reg __401719_401719;
   reg _401720_401720 ; 
   reg __401720_401720;
   reg _401721_401721 ; 
   reg __401721_401721;
   reg _401722_401722 ; 
   reg __401722_401722;
   reg _401723_401723 ; 
   reg __401723_401723;
   reg _401724_401724 ; 
   reg __401724_401724;
   reg _401725_401725 ; 
   reg __401725_401725;
   reg _401726_401726 ; 
   reg __401726_401726;
   reg _401727_401727 ; 
   reg __401727_401727;
   reg _401728_401728 ; 
   reg __401728_401728;
   reg _401729_401729 ; 
   reg __401729_401729;
   reg _401730_401730 ; 
   reg __401730_401730;
   reg _401731_401731 ; 
   reg __401731_401731;
   reg _401732_401732 ; 
   reg __401732_401732;
   reg _401733_401733 ; 
   reg __401733_401733;
   reg _401734_401734 ; 
   reg __401734_401734;
   reg _401735_401735 ; 
   reg __401735_401735;
   reg _401736_401736 ; 
   reg __401736_401736;
   reg _401737_401737 ; 
   reg __401737_401737;
   reg _401738_401738 ; 
   reg __401738_401738;
   reg _401739_401739 ; 
   reg __401739_401739;
   reg _401740_401740 ; 
   reg __401740_401740;
   reg _401741_401741 ; 
   reg __401741_401741;
   reg _401742_401742 ; 
   reg __401742_401742;
   reg _401743_401743 ; 
   reg __401743_401743;
   reg _401744_401744 ; 
   reg __401744_401744;
   reg _401745_401745 ; 
   reg __401745_401745;
   reg _401746_401746 ; 
   reg __401746_401746;
   reg _401747_401747 ; 
   reg __401747_401747;
   reg _401748_401748 ; 
   reg __401748_401748;
   reg _401749_401749 ; 
   reg __401749_401749;
   reg _401750_401750 ; 
   reg __401750_401750;
   reg _401751_401751 ; 
   reg __401751_401751;
   reg _401752_401752 ; 
   reg __401752_401752;
   reg _401753_401753 ; 
   reg __401753_401753;
   reg _401754_401754 ; 
   reg __401754_401754;
   reg _401755_401755 ; 
   reg __401755_401755;
   reg _401756_401756 ; 
   reg __401756_401756;
   reg _401757_401757 ; 
   reg __401757_401757;
   reg _401758_401758 ; 
   reg __401758_401758;
   reg _401759_401759 ; 
   reg __401759_401759;
   reg _401760_401760 ; 
   reg __401760_401760;
   reg _401761_401761 ; 
   reg __401761_401761;
   reg _401762_401762 ; 
   reg __401762_401762;
   reg _401763_401763 ; 
   reg __401763_401763;
   reg _401764_401764 ; 
   reg __401764_401764;
   reg _401765_401765 ; 
   reg __401765_401765;
   reg _401766_401766 ; 
   reg __401766_401766;
   reg _401767_401767 ; 
   reg __401767_401767;
   reg _401768_401768 ; 
   reg __401768_401768;
   reg _401769_401769 ; 
   reg __401769_401769;
   reg _401770_401770 ; 
   reg __401770_401770;
   reg _401771_401771 ; 
   reg __401771_401771;
   reg _401772_401772 ; 
   reg __401772_401772;
   reg _401773_401773 ; 
   reg __401773_401773;
   reg _401774_401774 ; 
   reg __401774_401774;
   reg _401775_401775 ; 
   reg __401775_401775;
   reg _401776_401776 ; 
   reg __401776_401776;
   reg _401777_401777 ; 
   reg __401777_401777;
   reg _401778_401778 ; 
   reg __401778_401778;
   reg _401779_401779 ; 
   reg __401779_401779;
   reg _401780_401780 ; 
   reg __401780_401780;
   reg _401781_401781 ; 
   reg __401781_401781;
   reg _401782_401782 ; 
   reg __401782_401782;
   reg _401783_401783 ; 
   reg __401783_401783;
   reg _401784_401784 ; 
   reg __401784_401784;
   reg _401785_401785 ; 
   reg __401785_401785;
   reg _401786_401786 ; 
   reg __401786_401786;
   reg _401787_401787 ; 
   reg __401787_401787;
   reg _401788_401788 ; 
   reg __401788_401788;
   reg _401789_401789 ; 
   reg __401789_401789;
   reg _401790_401790 ; 
   reg __401790_401790;
   reg _401791_401791 ; 
   reg __401791_401791;
   reg _401792_401792 ; 
   reg __401792_401792;
   reg _401793_401793 ; 
   reg __401793_401793;
   reg _401794_401794 ; 
   reg __401794_401794;
   reg _401795_401795 ; 
   reg __401795_401795;
   reg _401796_401796 ; 
   reg __401796_401796;
   reg _401797_401797 ; 
   reg __401797_401797;
   reg _401798_401798 ; 
   reg __401798_401798;
   reg _401799_401799 ; 
   reg __401799_401799;
   reg _401800_401800 ; 
   reg __401800_401800;
   reg _401801_401801 ; 
   reg __401801_401801;
   reg _401802_401802 ; 
   reg __401802_401802;
   reg _401803_401803 ; 
   reg __401803_401803;
   reg _401804_401804 ; 
   reg __401804_401804;
   reg _401805_401805 ; 
   reg __401805_401805;
   reg _401806_401806 ; 
   reg __401806_401806;
   reg _401807_401807 ; 
   reg __401807_401807;
   reg _401808_401808 ; 
   reg __401808_401808;
   reg _401809_401809 ; 
   reg __401809_401809;
   reg _401810_401810 ; 
   reg __401810_401810;
   reg _401811_401811 ; 
   reg __401811_401811;
   reg _401812_401812 ; 
   reg __401812_401812;
   reg _401813_401813 ; 
   reg __401813_401813;
   reg _401814_401814 ; 
   reg __401814_401814;
   reg _401815_401815 ; 
   reg __401815_401815;
   reg _401816_401816 ; 
   reg __401816_401816;
   reg _401817_401817 ; 
   reg __401817_401817;
   reg _401818_401818 ; 
   reg __401818_401818;
   reg _401819_401819 ; 
   reg __401819_401819;
   reg _401820_401820 ; 
   reg __401820_401820;
   reg _401821_401821 ; 
   reg __401821_401821;
   reg _401822_401822 ; 
   reg __401822_401822;
   reg _401823_401823 ; 
   reg __401823_401823;
   reg _401824_401824 ; 
   reg __401824_401824;
   reg _401825_401825 ; 
   reg __401825_401825;
   reg _401826_401826 ; 
   reg __401826_401826;
   reg _401827_401827 ; 
   reg __401827_401827;
   reg _401828_401828 ; 
   reg __401828_401828;
   reg _401829_401829 ; 
   reg __401829_401829;
   reg _401830_401830 ; 
   reg __401830_401830;
   reg _401831_401831 ; 
   reg __401831_401831;
   reg _401832_401832 ; 
   reg __401832_401832;
   reg _401833_401833 ; 
   reg __401833_401833;
   reg _401834_401834 ; 
   reg __401834_401834;
   reg _401835_401835 ; 
   reg __401835_401835;
   reg _401836_401836 ; 
   reg __401836_401836;
   reg _401837_401837 ; 
   reg __401837_401837;
   reg _401838_401838 ; 
   reg __401838_401838;
   reg _401839_401839 ; 
   reg __401839_401839;
   reg _401840_401840 ; 
   reg __401840_401840;
   reg _401841_401841 ; 
   reg __401841_401841;
   reg _401842_401842 ; 
   reg __401842_401842;
   reg _401843_401843 ; 
   reg __401843_401843;
   reg _401844_401844 ; 
   reg __401844_401844;
   reg _401845_401845 ; 
   reg __401845_401845;
   reg _401846_401846 ; 
   reg __401846_401846;
   reg _401847_401847 ; 
   reg __401847_401847;
   reg _401848_401848 ; 
   reg __401848_401848;
   reg _401849_401849 ; 
   reg __401849_401849;
   reg _401850_401850 ; 
   reg __401850_401850;
   reg _401851_401851 ; 
   reg __401851_401851;
   reg _401852_401852 ; 
   reg __401852_401852;
   reg _401853_401853 ; 
   reg __401853_401853;
   reg _401854_401854 ; 
   reg __401854_401854;
   reg _401855_401855 ; 
   reg __401855_401855;
   reg _401856_401856 ; 
   reg __401856_401856;
   reg _401857_401857 ; 
   reg __401857_401857;
   reg _401858_401858 ; 
   reg __401858_401858;
   reg _401859_401859 ; 
   reg __401859_401859;
   reg _401860_401860 ; 
   reg __401860_401860;
   reg _401861_401861 ; 
   reg __401861_401861;
   reg _401862_401862 ; 
   reg __401862_401862;
   reg _401863_401863 ; 
   reg __401863_401863;
   reg _401864_401864 ; 
   reg __401864_401864;
   reg _401865_401865 ; 
   reg __401865_401865;
   reg _401866_401866 ; 
   reg __401866_401866;
   reg _401867_401867 ; 
   reg __401867_401867;
   reg _401868_401868 ; 
   reg __401868_401868;
   reg _401869_401869 ; 
   reg __401869_401869;
   reg _401870_401870 ; 
   reg __401870_401870;
   reg _401871_401871 ; 
   reg __401871_401871;
   reg _401872_401872 ; 
   reg __401872_401872;
   reg _401873_401873 ; 
   reg __401873_401873;
   reg _401874_401874 ; 
   reg __401874_401874;
   reg _401875_401875 ; 
   reg __401875_401875;
   reg _401876_401876 ; 
   reg __401876_401876;
   reg _401877_401877 ; 
   reg __401877_401877;
   reg _401878_401878 ; 
   reg __401878_401878;
   reg _401879_401879 ; 
   reg __401879_401879;
   reg _401880_401880 ; 
   reg __401880_401880;
   reg _401881_401881 ; 
   reg __401881_401881;
   reg _401882_401882 ; 
   reg __401882_401882;
   reg _401883_401883 ; 
   reg __401883_401883;
   reg _401884_401884 ; 
   reg __401884_401884;
   reg _401885_401885 ; 
   reg __401885_401885;
   reg _401886_401886 ; 
   reg __401886_401886;
   reg _401887_401887 ; 
   reg __401887_401887;
   reg _401888_401888 ; 
   reg __401888_401888;
   reg _401889_401889 ; 
   reg __401889_401889;
   reg _401890_401890 ; 
   reg __401890_401890;
   reg _401891_401891 ; 
   reg __401891_401891;
   reg _401892_401892 ; 
   reg __401892_401892;
   reg _401893_401893 ; 
   reg __401893_401893;
   reg _401894_401894 ; 
   reg __401894_401894;
   reg _401895_401895 ; 
   reg __401895_401895;
   reg _401896_401896 ; 
   reg __401896_401896;
   reg _401897_401897 ; 
   reg __401897_401897;
   reg _401898_401898 ; 
   reg __401898_401898;
   reg _401899_401899 ; 
   reg __401899_401899;
   reg _401900_401900 ; 
   reg __401900_401900;
   reg _401901_401901 ; 
   reg __401901_401901;
   reg _401902_401902 ; 
   reg __401902_401902;
   reg _401903_401903 ; 
   reg __401903_401903;
   reg _401904_401904 ; 
   reg __401904_401904;
   reg _401905_401905 ; 
   reg __401905_401905;
   reg _401906_401906 ; 
   reg __401906_401906;
   reg _401907_401907 ; 
   reg __401907_401907;
   reg _401908_401908 ; 
   reg __401908_401908;
   reg _401909_401909 ; 
   reg __401909_401909;
   reg _401910_401910 ; 
   reg __401910_401910;
   reg _401911_401911 ; 
   reg __401911_401911;
   reg _401912_401912 ; 
   reg __401912_401912;
   reg _401913_401913 ; 
   reg __401913_401913;
   reg _401914_401914 ; 
   reg __401914_401914;
   reg _401915_401915 ; 
   reg __401915_401915;
   reg _401916_401916 ; 
   reg __401916_401916;
   reg _401917_401917 ; 
   reg __401917_401917;
   reg _401918_401918 ; 
   reg __401918_401918;
   reg _401919_401919 ; 
   reg __401919_401919;
   reg _401920_401920 ; 
   reg __401920_401920;
   reg _401921_401921 ; 
   reg __401921_401921;
   reg _401922_401922 ; 
   reg __401922_401922;
   reg _401923_401923 ; 
   reg __401923_401923;
   reg _401924_401924 ; 
   reg __401924_401924;
   reg _401925_401925 ; 
   reg __401925_401925;
   reg _401926_401926 ; 
   reg __401926_401926;
   reg _401927_401927 ; 
   reg __401927_401927;
   reg _401928_401928 ; 
   reg __401928_401928;
   reg _401929_401929 ; 
   reg __401929_401929;
   reg _401930_401930 ; 
   reg __401930_401930;
   reg _401931_401931 ; 
   reg __401931_401931;
   reg _401932_401932 ; 
   reg __401932_401932;
   reg _401933_401933 ; 
   reg __401933_401933;
   reg _401934_401934 ; 
   reg __401934_401934;
   reg _401935_401935 ; 
   reg __401935_401935;
   reg _401936_401936 ; 
   reg __401936_401936;
   reg _401937_401937 ; 
   reg __401937_401937;
   reg _401938_401938 ; 
   reg __401938_401938;
   reg _401939_401939 ; 
   reg __401939_401939;
   reg _401940_401940 ; 
   reg __401940_401940;
   reg _401941_401941 ; 
   reg __401941_401941;
   reg _401942_401942 ; 
   reg __401942_401942;
   reg _401943_401943 ; 
   reg __401943_401943;
   reg _401944_401944 ; 
   reg __401944_401944;
   reg _401945_401945 ; 
   reg __401945_401945;
   reg _401946_401946 ; 
   reg __401946_401946;
   reg _401947_401947 ; 
   reg __401947_401947;
   reg _401948_401948 ; 
   reg __401948_401948;
   reg _401949_401949 ; 
   reg __401949_401949;
   reg _401950_401950 ; 
   reg __401950_401950;
   reg _401951_401951 ; 
   reg __401951_401951;
   reg _401952_401952 ; 
   reg __401952_401952;
   reg _401953_401953 ; 
   reg __401953_401953;
   reg _401954_401954 ; 
   reg __401954_401954;
   reg _401955_401955 ; 
   reg __401955_401955;
   reg _401956_401956 ; 
   reg __401956_401956;
   reg _401957_401957 ; 
   reg __401957_401957;
   reg _401958_401958 ; 
   reg __401958_401958;
   reg _401959_401959 ; 
   reg __401959_401959;
   reg _401960_401960 ; 
   reg __401960_401960;
   reg _401961_401961 ; 
   reg __401961_401961;
   reg _401962_401962 ; 
   reg __401962_401962;
   reg _401963_401963 ; 
   reg __401963_401963;
   reg _401964_401964 ; 
   reg __401964_401964;
   reg _401965_401965 ; 
   reg __401965_401965;
   reg _401966_401966 ; 
   reg __401966_401966;
   reg _401967_401967 ; 
   reg __401967_401967;
   reg _401968_401968 ; 
   reg __401968_401968;
   reg _401969_401969 ; 
   reg __401969_401969;
   reg _401970_401970 ; 
   reg __401970_401970;
   reg _401971_401971 ; 
   reg __401971_401971;
   reg _401972_401972 ; 
   reg __401972_401972;
   reg _401973_401973 ; 
   reg __401973_401973;
   reg _401974_401974 ; 
   reg __401974_401974;
   reg _401975_401975 ; 
   reg __401975_401975;
   reg _401976_401976 ; 
   reg __401976_401976;
   reg _401977_401977 ; 
   reg __401977_401977;
   reg _401978_401978 ; 
   reg __401978_401978;
   reg _401979_401979 ; 
   reg __401979_401979;
   reg _401980_401980 ; 
   reg __401980_401980;
   reg _401981_401981 ; 
   reg __401981_401981;
   reg _401982_401982 ; 
   reg __401982_401982;
   reg _401983_401983 ; 
   reg __401983_401983;
   reg _401984_401984 ; 
   reg __401984_401984;
   reg _401985_401985 ; 
   reg __401985_401985;
   reg _401986_401986 ; 
   reg __401986_401986;
   reg _401987_401987 ; 
   reg __401987_401987;
   reg _401988_401988 ; 
   reg __401988_401988;
   reg _401989_401989 ; 
   reg __401989_401989;
   reg _401990_401990 ; 
   reg __401990_401990;
   reg _401991_401991 ; 
   reg __401991_401991;
   reg _401992_401992 ; 
   reg __401992_401992;
   reg _401993_401993 ; 
   reg __401993_401993;
   reg _401994_401994 ; 
   reg __401994_401994;
   reg _401995_401995 ; 
   reg __401995_401995;
   reg _401996_401996 ; 
   reg __401996_401996;
   reg _401997_401997 ; 
   reg __401997_401997;
   reg _401998_401998 ; 
   reg __401998_401998;
   reg _401999_401999 ; 
   reg __401999_401999;
   reg _402000_402000 ; 
   reg __402000_402000;
   reg _402001_402001 ; 
   reg __402001_402001;
   reg _402002_402002 ; 
   reg __402002_402002;
   reg _402003_402003 ; 
   reg __402003_402003;
   reg _402004_402004 ; 
   reg __402004_402004;
   reg _402005_402005 ; 
   reg __402005_402005;
   reg _402006_402006 ; 
   reg __402006_402006;
   reg _402007_402007 ; 
   reg __402007_402007;
   reg _402008_402008 ; 
   reg __402008_402008;
   reg _402009_402009 ; 
   reg __402009_402009;
   reg _402010_402010 ; 
   reg __402010_402010;
   reg _402011_402011 ; 
   reg __402011_402011;
   reg _402012_402012 ; 
   reg __402012_402012;
   reg _402013_402013 ; 
   reg __402013_402013;
   reg _402014_402014 ; 
   reg __402014_402014;
   reg _402015_402015 ; 
   reg __402015_402015;
   reg _402016_402016 ; 
   reg __402016_402016;
   reg _402017_402017 ; 
   reg __402017_402017;
   reg _402018_402018 ; 
   reg __402018_402018;
   reg _402019_402019 ; 
   reg __402019_402019;
   reg _402020_402020 ; 
   reg __402020_402020;
   reg _402021_402021 ; 
   reg __402021_402021;
   reg _402022_402022 ; 
   reg __402022_402022;
   reg _402023_402023 ; 
   reg __402023_402023;
   reg _402024_402024 ; 
   reg __402024_402024;
   reg _402025_402025 ; 
   reg __402025_402025;
   reg _402026_402026 ; 
   reg __402026_402026;
   reg _402027_402027 ; 
   reg __402027_402027;
   reg _402028_402028 ; 
   reg __402028_402028;
   reg _402029_402029 ; 
   reg __402029_402029;
   reg _402030_402030 ; 
   reg __402030_402030;
   reg _402031_402031 ; 
   reg __402031_402031;
   reg _402032_402032 ; 
   reg __402032_402032;
   reg _402033_402033 ; 
   reg __402033_402033;
   reg _402034_402034 ; 
   reg __402034_402034;
   reg _402035_402035 ; 
   reg __402035_402035;
   reg _402036_402036 ; 
   reg __402036_402036;
   reg _402037_402037 ; 
   reg __402037_402037;
   reg _402038_402038 ; 
   reg __402038_402038;
   reg _402039_402039 ; 
   reg __402039_402039;
   reg _402040_402040 ; 
   reg __402040_402040;
   reg _402041_402041 ; 
   reg __402041_402041;
   reg _402042_402042 ; 
   reg __402042_402042;
   reg _402043_402043 ; 
   reg __402043_402043;
   reg _402044_402044 ; 
   reg __402044_402044;
   reg _402045_402045 ; 
   reg __402045_402045;
   reg _402046_402046 ; 
   reg __402046_402046;
   reg _402047_402047 ; 
   reg __402047_402047;
   reg _402048_402048 ; 
   reg __402048_402048;
   reg _402049_402049 ; 
   reg __402049_402049;
   reg _402050_402050 ; 
   reg __402050_402050;
   reg _402051_402051 ; 
   reg __402051_402051;
   reg _402052_402052 ; 
   reg __402052_402052;
   reg _402053_402053 ; 
   reg __402053_402053;
   reg _402054_402054 ; 
   reg __402054_402054;
   reg _402055_402055 ; 
   reg __402055_402055;
   reg _402056_402056 ; 
   reg __402056_402056;
   reg _402057_402057 ; 
   reg __402057_402057;
   reg _402058_402058 ; 
   reg __402058_402058;
   reg _402059_402059 ; 
   reg __402059_402059;
   reg _402060_402060 ; 
   reg __402060_402060;
   reg _402061_402061 ; 
   reg __402061_402061;
   reg _402062_402062 ; 
   reg __402062_402062;
   reg _402063_402063 ; 
   reg __402063_402063;
   reg _402064_402064 ; 
   reg __402064_402064;
   reg _402065_402065 ; 
   reg __402065_402065;
   reg _402066_402066 ; 
   reg __402066_402066;
   reg _402067_402067 ; 
   reg __402067_402067;
   reg _402068_402068 ; 
   reg __402068_402068;
   reg _402069_402069 ; 
   reg __402069_402069;
   reg _402070_402070 ; 
   reg __402070_402070;
   reg _402071_402071 ; 
   reg __402071_402071;
   reg _402072_402072 ; 
   reg __402072_402072;
   reg _402073_402073 ; 
   reg __402073_402073;
   reg _402074_402074 ; 
   reg __402074_402074;
   reg _402075_402075 ; 
   reg __402075_402075;
   reg _402076_402076 ; 
   reg __402076_402076;
   reg _402077_402077 ; 
   reg __402077_402077;
   reg _402078_402078 ; 
   reg __402078_402078;
   reg _402079_402079 ; 
   reg __402079_402079;
   reg _402080_402080 ; 
   reg __402080_402080;
   reg _402081_402081 ; 
   reg __402081_402081;
   reg _402082_402082 ; 
   reg __402082_402082;
   reg _402083_402083 ; 
   reg __402083_402083;
   reg _402084_402084 ; 
   reg __402084_402084;
   reg _402085_402085 ; 
   reg __402085_402085;
   reg _402086_402086 ; 
   reg __402086_402086;
   reg _402087_402087 ; 
   reg __402087_402087;
   reg _402088_402088 ; 
   reg __402088_402088;
   reg _402089_402089 ; 
   reg __402089_402089;
   reg _402090_402090 ; 
   reg __402090_402090;
   reg _402091_402091 ; 
   reg __402091_402091;
   reg _402092_402092 ; 
   reg __402092_402092;
   reg _402093_402093 ; 
   reg __402093_402093;
   reg _402094_402094 ; 
   reg __402094_402094;
   reg _402095_402095 ; 
   reg __402095_402095;
   reg _402096_402096 ; 
   reg __402096_402096;
   reg _402097_402097 ; 
   reg __402097_402097;
   reg _402098_402098 ; 
   reg __402098_402098;
   reg _402099_402099 ; 
   reg __402099_402099;
   reg _402100_402100 ; 
   reg __402100_402100;
   reg _402101_402101 ; 
   reg __402101_402101;
   reg _402102_402102 ; 
   reg __402102_402102;
   reg _402103_402103 ; 
   reg __402103_402103;
   reg _402104_402104 ; 
   reg __402104_402104;
   reg _402105_402105 ; 
   reg __402105_402105;
   reg _402106_402106 ; 
   reg __402106_402106;
   reg _402107_402107 ; 
   reg __402107_402107;
   reg _402108_402108 ; 
   reg __402108_402108;
   reg _402109_402109 ; 
   reg __402109_402109;
   reg _402110_402110 ; 
   reg __402110_402110;
   reg _402111_402111 ; 
   reg __402111_402111;
   reg _402112_402112 ; 
   reg __402112_402112;
   reg _402113_402113 ; 
   reg __402113_402113;
   reg _402114_402114 ; 
   reg __402114_402114;
   reg _402115_402115 ; 
   reg __402115_402115;
   reg _402116_402116 ; 
   reg __402116_402116;
   reg _402117_402117 ; 
   reg __402117_402117;
   reg _402118_402118 ; 
   reg __402118_402118;
   reg _402119_402119 ; 
   reg __402119_402119;
   reg _402120_402120 ; 
   reg __402120_402120;
   reg _402121_402121 ; 
   reg __402121_402121;
   reg _402122_402122 ; 
   reg __402122_402122;
   reg _402123_402123 ; 
   reg __402123_402123;
   reg _402124_402124 ; 
   reg __402124_402124;
   reg _402125_402125 ; 
   reg __402125_402125;
   reg _402126_402126 ; 
   reg __402126_402126;
   reg _402127_402127 ; 
   reg __402127_402127;
   reg _402128_402128 ; 
   reg __402128_402128;
   reg _402129_402129 ; 
   reg __402129_402129;
   reg _402130_402130 ; 
   reg __402130_402130;
   reg _402131_402131 ; 
   reg __402131_402131;
   reg _402132_402132 ; 
   reg __402132_402132;
   reg _402133_402133 ; 
   reg __402133_402133;
   reg _402134_402134 ; 
   reg __402134_402134;
   reg _402135_402135 ; 
   reg __402135_402135;
   reg _402136_402136 ; 
   reg __402136_402136;
   reg _402137_402137 ; 
   reg __402137_402137;
   reg _402138_402138 ; 
   reg __402138_402138;
   reg _402139_402139 ; 
   reg __402139_402139;
   reg _402140_402140 ; 
   reg __402140_402140;
   reg _402141_402141 ; 
   reg __402141_402141;
   reg _402142_402142 ; 
   reg __402142_402142;
   reg _402143_402143 ; 
   reg __402143_402143;
   reg _402144_402144 ; 
   reg __402144_402144;
   reg _402145_402145 ; 
   reg __402145_402145;
   reg _402146_402146 ; 
   reg __402146_402146;
   reg _402147_402147 ; 
   reg __402147_402147;
   reg _402148_402148 ; 
   reg __402148_402148;
   reg _402149_402149 ; 
   reg __402149_402149;
   reg _402150_402150 ; 
   reg __402150_402150;
   reg _402151_402151 ; 
   reg __402151_402151;
   reg _402152_402152 ; 
   reg __402152_402152;
   reg _402153_402153 ; 
   reg __402153_402153;
   reg _402154_402154 ; 
   reg __402154_402154;
   reg _402155_402155 ; 
   reg __402155_402155;
   reg _402156_402156 ; 
   reg __402156_402156;
   reg _402157_402157 ; 
   reg __402157_402157;
   reg _402158_402158 ; 
   reg __402158_402158;
   reg _402159_402159 ; 
   reg __402159_402159;
   reg _402160_402160 ; 
   reg __402160_402160;
   reg _402161_402161 ; 
   reg __402161_402161;
   reg _402162_402162 ; 
   reg __402162_402162;
   reg _402163_402163 ; 
   reg __402163_402163;
   reg _402164_402164 ; 
   reg __402164_402164;
   reg _402165_402165 ; 
   reg __402165_402165;
   reg _402166_402166 ; 
   reg __402166_402166;
   reg _402167_402167 ; 
   reg __402167_402167;
   reg _402168_402168 ; 
   reg __402168_402168;
   reg _402169_402169 ; 
   reg __402169_402169;
   reg _402170_402170 ; 
   reg __402170_402170;
   reg _402171_402171 ; 
   reg __402171_402171;
   reg _402172_402172 ; 
   reg __402172_402172;
   reg _402173_402173 ; 
   reg __402173_402173;
   reg _402174_402174 ; 
   reg __402174_402174;
   reg _402175_402175 ; 
   reg __402175_402175;
   reg _402176_402176 ; 
   reg __402176_402176;
   reg _402177_402177 ; 
   reg __402177_402177;
   reg _402178_402178 ; 
   reg __402178_402178;
   reg _402179_402179 ; 
   reg __402179_402179;
   reg _402180_402180 ; 
   reg __402180_402180;
   reg _402181_402181 ; 
   reg __402181_402181;
   reg _402182_402182 ; 
   reg __402182_402182;
   reg _402183_402183 ; 
   reg __402183_402183;
   reg _402184_402184 ; 
   reg __402184_402184;
   reg _402185_402185 ; 
   reg __402185_402185;
   reg _402186_402186 ; 
   reg __402186_402186;
   reg _402187_402187 ; 
   reg __402187_402187;
   reg _402188_402188 ; 
   reg __402188_402188;
   reg _402189_402189 ; 
   reg __402189_402189;
   reg _402190_402190 ; 
   reg __402190_402190;
   reg _402191_402191 ; 
   reg __402191_402191;
   reg _402192_402192 ; 
   reg __402192_402192;
   reg _402193_402193 ; 
   reg __402193_402193;
   reg _402194_402194 ; 
   reg __402194_402194;
   reg _402195_402195 ; 
   reg __402195_402195;
   reg _402196_402196 ; 
   reg __402196_402196;
   reg _402197_402197 ; 
   reg __402197_402197;
   reg _402198_402198 ; 
   reg __402198_402198;
   reg _402199_402199 ; 
   reg __402199_402199;
   reg _402200_402200 ; 
   reg __402200_402200;
   reg _402201_402201 ; 
   reg __402201_402201;
   reg _402202_402202 ; 
   reg __402202_402202;
   reg _402203_402203 ; 
   reg __402203_402203;
   reg _402204_402204 ; 
   reg __402204_402204;
   reg _402205_402205 ; 
   reg __402205_402205;
   reg _402206_402206 ; 
   reg __402206_402206;
   reg _402207_402207 ; 
   reg __402207_402207;
   reg _402208_402208 ; 
   reg __402208_402208;
   reg _402209_402209 ; 
   reg __402209_402209;
   reg _402210_402210 ; 
   reg __402210_402210;
   reg _402211_402211 ; 
   reg __402211_402211;
   reg _402212_402212 ; 
   reg __402212_402212;
   reg _402213_402213 ; 
   reg __402213_402213;
   reg _402214_402214 ; 
   reg __402214_402214;
   reg _402215_402215 ; 
   reg __402215_402215;
   reg _402216_402216 ; 
   reg __402216_402216;
   reg _402217_402217 ; 
   reg __402217_402217;
   reg _402218_402218 ; 
   reg __402218_402218;
   reg _402219_402219 ; 
   reg __402219_402219;
   reg _402220_402220 ; 
   reg __402220_402220;
   reg _402221_402221 ; 
   reg __402221_402221;
   reg _402222_402222 ; 
   reg __402222_402222;
   reg _402223_402223 ; 
   reg __402223_402223;
   reg _402224_402224 ; 
   reg __402224_402224;
   reg _402225_402225 ; 
   reg __402225_402225;
   reg _402226_402226 ; 
   reg __402226_402226;
   reg _402227_402227 ; 
   reg __402227_402227;
   reg _402228_402228 ; 
   reg __402228_402228;
   reg _402229_402229 ; 
   reg __402229_402229;
   reg _402230_402230 ; 
   reg __402230_402230;
   reg _402231_402231 ; 
   reg __402231_402231;
   reg _402232_402232 ; 
   reg __402232_402232;
   reg _402233_402233 ; 
   reg __402233_402233;
   reg _402234_402234 ; 
   reg __402234_402234;
   reg _402235_402235 ; 
   reg __402235_402235;
   reg _402236_402236 ; 
   reg __402236_402236;
   reg _402237_402237 ; 
   reg __402237_402237;
   reg _402238_402238 ; 
   reg __402238_402238;
   reg _402239_402239 ; 
   reg __402239_402239;
   reg _402240_402240 ; 
   reg __402240_402240;
   reg _402241_402241 ; 
   reg __402241_402241;
   reg _402242_402242 ; 
   reg __402242_402242;
   reg _402243_402243 ; 
   reg __402243_402243;
   reg _402244_402244 ; 
   reg __402244_402244;
   reg _402245_402245 ; 
   reg __402245_402245;
   reg _402246_402246 ; 
   reg __402246_402246;
   reg _402247_402247 ; 
   reg __402247_402247;
   reg _402248_402248 ; 
   reg __402248_402248;
   reg _402249_402249 ; 
   reg __402249_402249;
   reg _402250_402250 ; 
   reg __402250_402250;
   reg _402251_402251 ; 
   reg __402251_402251;
   reg _402252_402252 ; 
   reg __402252_402252;
   reg _402253_402253 ; 
   reg __402253_402253;
   reg _402254_402254 ; 
   reg __402254_402254;
   reg _402255_402255 ; 
   reg __402255_402255;
   reg _402256_402256 ; 
   reg __402256_402256;
   reg _402257_402257 ; 
   reg __402257_402257;
   reg _402258_402258 ; 
   reg __402258_402258;
   reg _402259_402259 ; 
   reg __402259_402259;
   reg _402260_402260 ; 
   reg __402260_402260;
   reg _402261_402261 ; 
   reg __402261_402261;
   reg _402262_402262 ; 
   reg __402262_402262;
   reg _402263_402263 ; 
   reg __402263_402263;
   reg _402264_402264 ; 
   reg __402264_402264;
   reg _402265_402265 ; 
   reg __402265_402265;
   reg _402266_402266 ; 
   reg __402266_402266;
   reg _402267_402267 ; 
   reg __402267_402267;
   reg _402268_402268 ; 
   reg __402268_402268;
   reg _402269_402269 ; 
   reg __402269_402269;
   reg _402270_402270 ; 
   reg __402270_402270;
   reg _402271_402271 ; 
   reg __402271_402271;
   reg _402272_402272 ; 
   reg __402272_402272;
   reg _402273_402273 ; 
   reg __402273_402273;
   reg _402274_402274 ; 
   reg __402274_402274;
   reg _402275_402275 ; 
   reg __402275_402275;
   reg _402276_402276 ; 
   reg __402276_402276;
   reg _402277_402277 ; 
   reg __402277_402277;
   reg _402278_402278 ; 
   reg __402278_402278;
   reg _402279_402279 ; 
   reg __402279_402279;
   reg _402280_402280 ; 
   reg __402280_402280;
   reg _402281_402281 ; 
   reg __402281_402281;
   reg _402282_402282 ; 
   reg __402282_402282;
   reg _402283_402283 ; 
   reg __402283_402283;
   reg _402284_402284 ; 
   reg __402284_402284;
   reg _402285_402285 ; 
   reg __402285_402285;
   reg _402286_402286 ; 
   reg __402286_402286;
   reg _402287_402287 ; 
   reg __402287_402287;
   reg _402288_402288 ; 
   reg __402288_402288;
   reg _402289_402289 ; 
   reg __402289_402289;
   reg _402290_402290 ; 
   reg __402290_402290;
   reg _402291_402291 ; 
   reg __402291_402291;
   reg _402292_402292 ; 
   reg __402292_402292;
   reg _402293_402293 ; 
   reg __402293_402293;
   reg _402294_402294 ; 
   reg __402294_402294;
   reg _402295_402295 ; 
   reg __402295_402295;
   reg _402296_402296 ; 
   reg __402296_402296;
   reg _402297_402297 ; 
   reg __402297_402297;
   reg _402298_402298 ; 
   reg __402298_402298;
   reg _402299_402299 ; 
   reg __402299_402299;
   reg _402300_402300 ; 
   reg __402300_402300;
   reg _402301_402301 ; 
   reg __402301_402301;
   reg _402302_402302 ; 
   reg __402302_402302;
   reg _402303_402303 ; 
   reg __402303_402303;
   reg _402304_402304 ; 
   reg __402304_402304;
   reg _402305_402305 ; 
   reg __402305_402305;
   reg _402306_402306 ; 
   reg __402306_402306;
   reg _402307_402307 ; 
   reg __402307_402307;
   reg _402308_402308 ; 
   reg __402308_402308;
   reg _402309_402309 ; 
   reg __402309_402309;
   reg _402310_402310 ; 
   reg __402310_402310;
   reg _402311_402311 ; 
   reg __402311_402311;
   reg _402312_402312 ; 
   reg __402312_402312;
   reg _402313_402313 ; 
   reg __402313_402313;
   reg _402314_402314 ; 
   reg __402314_402314;
   reg _402315_402315 ; 
   reg __402315_402315;
   reg _402316_402316 ; 
   reg __402316_402316;
   reg _402317_402317 ; 
   reg __402317_402317;
   reg _402318_402318 ; 
   reg __402318_402318;
   reg _402319_402319 ; 
   reg __402319_402319;
   reg _402320_402320 ; 
   reg __402320_402320;
   reg _402321_402321 ; 
   reg __402321_402321;
   reg _402322_402322 ; 
   reg __402322_402322;
   reg _402323_402323 ; 
   reg __402323_402323;
   reg _402324_402324 ; 
   reg __402324_402324;
   reg _402325_402325 ; 
   reg __402325_402325;
   reg _402326_402326 ; 
   reg __402326_402326;
   reg _402327_402327 ; 
   reg __402327_402327;
   reg _402328_402328 ; 
   reg __402328_402328;
   reg _402329_402329 ; 
   reg __402329_402329;
   reg _402330_402330 ; 
   reg __402330_402330;
   reg _402331_402331 ; 
   reg __402331_402331;
   reg _402332_402332 ; 
   reg __402332_402332;
   reg _402333_402333 ; 
   reg __402333_402333;
   reg _402334_402334 ; 
   reg __402334_402334;
   reg _402335_402335 ; 
   reg __402335_402335;
   reg _402336_402336 ; 
   reg __402336_402336;
   reg _402337_402337 ; 
   reg __402337_402337;
   reg _402338_402338 ; 
   reg __402338_402338;
   reg _402339_402339 ; 
   reg __402339_402339;
   reg _402340_402340 ; 
   reg __402340_402340;
   reg _402341_402341 ; 
   reg __402341_402341;
   reg _402342_402342 ; 
   reg __402342_402342;
   reg _402343_402343 ; 
   reg __402343_402343;
   reg _402344_402344 ; 
   reg __402344_402344;
   reg _402345_402345 ; 
   reg __402345_402345;
   reg _402346_402346 ; 
   reg __402346_402346;
   reg _402347_402347 ; 
   reg __402347_402347;
   reg _402348_402348 ; 
   reg __402348_402348;
   reg _402349_402349 ; 
   reg __402349_402349;
   reg _402350_402350 ; 
   reg __402350_402350;
   reg _402351_402351 ; 
   reg __402351_402351;
   reg _402352_402352 ; 
   reg __402352_402352;
   reg _402353_402353 ; 
   reg __402353_402353;
   reg _402354_402354 ; 
   reg __402354_402354;
   reg _402355_402355 ; 
   reg __402355_402355;
   reg _402356_402356 ; 
   reg __402356_402356;
   reg _402357_402357 ; 
   reg __402357_402357;
   reg _402358_402358 ; 
   reg __402358_402358;
   reg _402359_402359 ; 
   reg __402359_402359;
   reg _402360_402360 ; 
   reg __402360_402360;
   reg _402361_402361 ; 
   reg __402361_402361;
   reg _402362_402362 ; 
   reg __402362_402362;
   reg _402363_402363 ; 
   reg __402363_402363;
   reg _402364_402364 ; 
   reg __402364_402364;
   reg _402365_402365 ; 
   reg __402365_402365;
   reg _402366_402366 ; 
   reg __402366_402366;
   reg _402367_402367 ; 
   reg __402367_402367;
   reg _402368_402368 ; 
   reg __402368_402368;
   reg _402369_402369 ; 
   reg __402369_402369;
   reg _402370_402370 ; 
   reg __402370_402370;
   reg _402371_402371 ; 
   reg __402371_402371;
   reg _402372_402372 ; 
   reg __402372_402372;
   reg _402373_402373 ; 
   reg __402373_402373;
   reg _402374_402374 ; 
   reg __402374_402374;
   reg _402375_402375 ; 
   reg __402375_402375;
   reg _402376_402376 ; 
   reg __402376_402376;
   reg _402377_402377 ; 
   reg __402377_402377;
   reg _402378_402378 ; 
   reg __402378_402378;
   reg _402379_402379 ; 
   reg __402379_402379;
   reg _402380_402380 ; 
   reg __402380_402380;
   reg _402381_402381 ; 
   reg __402381_402381;
   reg _402382_402382 ; 
   reg __402382_402382;
   reg _402383_402383 ; 
   reg __402383_402383;
   reg _402384_402384 ; 
   reg __402384_402384;
   reg _402385_402385 ; 
   reg __402385_402385;
   reg _402386_402386 ; 
   reg __402386_402386;
   reg _402387_402387 ; 
   reg __402387_402387;
   reg _402388_402388 ; 
   reg __402388_402388;
   reg _402389_402389 ; 
   reg __402389_402389;
   reg _402390_402390 ; 
   reg __402390_402390;
   reg _402391_402391 ; 
   reg __402391_402391;
   reg _402392_402392 ; 
   reg __402392_402392;
   reg _402393_402393 ; 
   reg __402393_402393;
   reg _402394_402394 ; 
   reg __402394_402394;
   reg _402395_402395 ; 
   reg __402395_402395;
   reg _402396_402396 ; 
   reg __402396_402396;
   reg _402397_402397 ; 
   reg __402397_402397;
   reg _402398_402398 ; 
   reg __402398_402398;
   reg _402399_402399 ; 
   reg __402399_402399;
   reg _402400_402400 ; 
   reg __402400_402400;
   reg _402401_402401 ; 
   reg __402401_402401;
   reg _402402_402402 ; 
   reg __402402_402402;
   reg _402403_402403 ; 
   reg __402403_402403;
   reg _402404_402404 ; 
   reg __402404_402404;
   reg _402405_402405 ; 
   reg __402405_402405;
   reg _402406_402406 ; 
   reg __402406_402406;
   reg _402407_402407 ; 
   reg __402407_402407;
   reg _402408_402408 ; 
   reg __402408_402408;
   reg _402409_402409 ; 
   reg __402409_402409;
   reg _402410_402410 ; 
   reg __402410_402410;
   reg _402411_402411 ; 
   reg __402411_402411;
   reg _402412_402412 ; 
   reg __402412_402412;
   reg _402413_402413 ; 
   reg __402413_402413;
   reg _402414_402414 ; 
   reg __402414_402414;
   reg _402415_402415 ; 
   reg __402415_402415;
   reg _402416_402416 ; 
   reg __402416_402416;
   reg _402417_402417 ; 
   reg __402417_402417;
   reg _402418_402418 ; 
   reg __402418_402418;
   reg _402419_402419 ; 
   reg __402419_402419;
   reg _402420_402420 ; 
   reg __402420_402420;
   reg _402421_402421 ; 
   reg __402421_402421;
   reg _402422_402422 ; 
   reg __402422_402422;
   reg _402423_402423 ; 
   reg __402423_402423;
   reg _402424_402424 ; 
   reg __402424_402424;
   reg _402425_402425 ; 
   reg __402425_402425;
   reg _402426_402426 ; 
   reg __402426_402426;
   reg _402427_402427 ; 
   reg __402427_402427;
   reg _402428_402428 ; 
   reg __402428_402428;
   reg _402429_402429 ; 
   reg __402429_402429;
   reg _402430_402430 ; 
   reg __402430_402430;
   reg _402431_402431 ; 
   reg __402431_402431;
   reg _402432_402432 ; 
   reg __402432_402432;
   reg _402433_402433 ; 
   reg __402433_402433;
   reg _402434_402434 ; 
   reg __402434_402434;
   reg _402435_402435 ; 
   reg __402435_402435;
   reg _402436_402436 ; 
   reg __402436_402436;
   reg _402437_402437 ; 
   reg __402437_402437;
   reg _402438_402438 ; 
   reg __402438_402438;
   reg _402439_402439 ; 
   reg __402439_402439;
   reg _402440_402440 ; 
   reg __402440_402440;
   reg _402441_402441 ; 
   reg __402441_402441;
   reg _402442_402442 ; 
   reg __402442_402442;
   reg _402443_402443 ; 
   reg __402443_402443;
   reg _402444_402444 ; 
   reg __402444_402444;
   reg _402445_402445 ; 
   reg __402445_402445;
   reg _402446_402446 ; 
   reg __402446_402446;
   reg _402447_402447 ; 
   reg __402447_402447;
   reg _402448_402448 ; 
   reg __402448_402448;
   reg _402449_402449 ; 
   reg __402449_402449;
   reg _402450_402450 ; 
   reg __402450_402450;
   reg _402451_402451 ; 
   reg __402451_402451;
   reg _402452_402452 ; 
   reg __402452_402452;
   reg _402453_402453 ; 
   reg __402453_402453;
   reg _402454_402454 ; 
   reg __402454_402454;
   reg _402455_402455 ; 
   reg __402455_402455;
   reg _402456_402456 ; 
   reg __402456_402456;
   reg _402457_402457 ; 
   reg __402457_402457;
   reg _402458_402458 ; 
   reg __402458_402458;
   reg _402459_402459 ; 
   reg __402459_402459;
   reg _402460_402460 ; 
   reg __402460_402460;
   reg _402461_402461 ; 
   reg __402461_402461;
   reg _402462_402462 ; 
   reg __402462_402462;
   reg _402463_402463 ; 
   reg __402463_402463;
   reg _402464_402464 ; 
   reg __402464_402464;
   reg _402465_402465 ; 
   reg __402465_402465;
   reg _402466_402466 ; 
   reg __402466_402466;
   reg _402467_402467 ; 
   reg __402467_402467;
   reg _402468_402468 ; 
   reg __402468_402468;
   reg _402469_402469 ; 
   reg __402469_402469;
   reg _402470_402470 ; 
   reg __402470_402470;
   reg _402471_402471 ; 
   reg __402471_402471;
   reg _402472_402472 ; 
   reg __402472_402472;
   reg _402473_402473 ; 
   reg __402473_402473;
   reg _402474_402474 ; 
   reg __402474_402474;
   reg _402475_402475 ; 
   reg __402475_402475;
   reg _402476_402476 ; 
   reg __402476_402476;
   reg _402477_402477 ; 
   reg __402477_402477;
   reg _402478_402478 ; 
   reg __402478_402478;
   reg _402479_402479 ; 
   reg __402479_402479;
   reg _402480_402480 ; 
   reg __402480_402480;
   reg _402481_402481 ; 
   reg __402481_402481;
   reg _402482_402482 ; 
   reg __402482_402482;
   reg _402483_402483 ; 
   reg __402483_402483;
   reg _402484_402484 ; 
   reg __402484_402484;
   reg _402485_402485 ; 
   reg __402485_402485;
   reg _402486_402486 ; 
   reg __402486_402486;
   reg _402487_402487 ; 
   reg __402487_402487;
   reg _402488_402488 ; 
   reg __402488_402488;
   reg _402489_402489 ; 
   reg __402489_402489;
   reg _402490_402490 ; 
   reg __402490_402490;
   reg _402491_402491 ; 
   reg __402491_402491;
   reg _402492_402492 ; 
   reg __402492_402492;
   reg _402493_402493 ; 
   reg __402493_402493;
   reg _402494_402494 ; 
   reg __402494_402494;
   reg _402495_402495 ; 
   reg __402495_402495;
   reg _402496_402496 ; 
   reg __402496_402496;
   reg _402497_402497 ; 
   reg __402497_402497;
   reg _402498_402498 ; 
   reg __402498_402498;
   reg _402499_402499 ; 
   reg __402499_402499;
   reg _402500_402500 ; 
   reg __402500_402500;
   reg _402501_402501 ; 
   reg __402501_402501;
   reg _402502_402502 ; 
   reg __402502_402502;
   reg _402503_402503 ; 
   reg __402503_402503;
   reg _402504_402504 ; 
   reg __402504_402504;
   reg _402505_402505 ; 
   reg __402505_402505;
   reg _402506_402506 ; 
   reg __402506_402506;
   reg _402507_402507 ; 
   reg __402507_402507;
   reg _402508_402508 ; 
   reg __402508_402508;
   reg _402509_402509 ; 
   reg __402509_402509;
   reg _402510_402510 ; 
   reg __402510_402510;
   reg _402511_402511 ; 
   reg __402511_402511;
   reg _402512_402512 ; 
   reg __402512_402512;
   reg _402513_402513 ; 
   reg __402513_402513;
   reg _402514_402514 ; 
   reg __402514_402514;
   reg _402515_402515 ; 
   reg __402515_402515;
   reg _402516_402516 ; 
   reg __402516_402516;
   reg _402517_402517 ; 
   reg __402517_402517;
   reg _402518_402518 ; 
   reg __402518_402518;
   reg _402519_402519 ; 
   reg __402519_402519;
   reg _402520_402520 ; 
   reg __402520_402520;
   reg _402521_402521 ; 
   reg __402521_402521;
   reg _402522_402522 ; 
   reg __402522_402522;
   reg _402523_402523 ; 
   reg __402523_402523;
   reg _402524_402524 ; 
   reg __402524_402524;
   reg _402525_402525 ; 
   reg __402525_402525;
   reg _402526_402526 ; 
   reg __402526_402526;
   reg _402527_402527 ; 
   reg __402527_402527;
   reg _402528_402528 ; 
   reg __402528_402528;
   reg _402529_402529 ; 
   reg __402529_402529;
   reg _402530_402530 ; 
   reg __402530_402530;
   reg _402531_402531 ; 
   reg __402531_402531;
   reg _402532_402532 ; 
   reg __402532_402532;
   reg _402533_402533 ; 
   reg __402533_402533;
   reg _402534_402534 ; 
   reg __402534_402534;
   reg _402535_402535 ; 
   reg __402535_402535;
   reg _402536_402536 ; 
   reg __402536_402536;
   reg _402537_402537 ; 
   reg __402537_402537;
   reg _402538_402538 ; 
   reg __402538_402538;
   reg _402539_402539 ; 
   reg __402539_402539;
   reg _402540_402540 ; 
   reg __402540_402540;
   reg _402541_402541 ; 
   reg __402541_402541;
   reg _402542_402542 ; 
   reg __402542_402542;
   reg _402543_402543 ; 
   reg __402543_402543;
   reg _402544_402544 ; 
   reg __402544_402544;
   reg _402545_402545 ; 
   reg __402545_402545;
   reg _402546_402546 ; 
   reg __402546_402546;
   reg _402547_402547 ; 
   reg __402547_402547;
   reg _402548_402548 ; 
   reg __402548_402548;
   reg _402549_402549 ; 
   reg __402549_402549;
   reg _402550_402550 ; 
   reg __402550_402550;
   reg _402551_402551 ; 
   reg __402551_402551;
   reg _402552_402552 ; 
   reg __402552_402552;
   reg _402553_402553 ; 
   reg __402553_402553;
   reg _402554_402554 ; 
   reg __402554_402554;
   reg _402555_402555 ; 
   reg __402555_402555;
   reg _402556_402556 ; 
   reg __402556_402556;
   reg _402557_402557 ; 
   reg __402557_402557;
   reg _402558_402558 ; 
   reg __402558_402558;
   reg _402559_402559 ; 
   reg __402559_402559;
   reg _402560_402560 ; 
   reg __402560_402560;
   reg _402561_402561 ; 
   reg __402561_402561;
   reg _402562_402562 ; 
   reg __402562_402562;
   reg _402563_402563 ; 
   reg __402563_402563;
   reg _402564_402564 ; 
   reg __402564_402564;
   reg _402565_402565 ; 
   reg __402565_402565;
   reg _402566_402566 ; 
   reg __402566_402566;
   reg _402567_402567 ; 
   reg __402567_402567;
   reg _402568_402568 ; 
   reg __402568_402568;
   reg _402569_402569 ; 
   reg __402569_402569;
   reg _402570_402570 ; 
   reg __402570_402570;
   reg _402571_402571 ; 
   reg __402571_402571;
   reg _402572_402572 ; 
   reg __402572_402572;
   reg _402573_402573 ; 
   reg __402573_402573;
   reg _402574_402574 ; 
   reg __402574_402574;
   reg _402575_402575 ; 
   reg __402575_402575;
   reg _402576_402576 ; 
   reg __402576_402576;
   reg _402577_402577 ; 
   reg __402577_402577;
   reg _402578_402578 ; 
   reg __402578_402578;
   reg _402579_402579 ; 
   reg __402579_402579;
   reg _402580_402580 ; 
   reg __402580_402580;
   reg _402581_402581 ; 
   reg __402581_402581;
   reg _402582_402582 ; 
   reg __402582_402582;
   reg _402583_402583 ; 
   reg __402583_402583;
   reg _402584_402584 ; 
   reg __402584_402584;
   reg _402585_402585 ; 
   reg __402585_402585;
   reg _402586_402586 ; 
   reg __402586_402586;
   reg _402587_402587 ; 
   reg __402587_402587;
   reg _402588_402588 ; 
   reg __402588_402588;
   reg _402589_402589 ; 
   reg __402589_402589;
   reg _402590_402590 ; 
   reg __402590_402590;
   reg _402591_402591 ; 
   reg __402591_402591;
   reg _402592_402592 ; 
   reg __402592_402592;
   reg _402593_402593 ; 
   reg __402593_402593;
   reg _402594_402594 ; 
   reg __402594_402594;
   reg _402595_402595 ; 
   reg __402595_402595;
   reg _402596_402596 ; 
   reg __402596_402596;
   reg _402597_402597 ; 
   reg __402597_402597;
   reg _402598_402598 ; 
   reg __402598_402598;
   reg _402599_402599 ; 
   reg __402599_402599;
   reg _402600_402600 ; 
   reg __402600_402600;
   reg _402601_402601 ; 
   reg __402601_402601;
   reg _402602_402602 ; 
   reg __402602_402602;
   reg _402603_402603 ; 
   reg __402603_402603;
   reg _402604_402604 ; 
   reg __402604_402604;
   reg _402605_402605 ; 
   reg __402605_402605;
   reg _402606_402606 ; 
   reg __402606_402606;
   reg _402607_402607 ; 
   reg __402607_402607;
   reg _402608_402608 ; 
   reg __402608_402608;
   reg _402609_402609 ; 
   reg __402609_402609;
   reg _402610_402610 ; 
   reg __402610_402610;
   reg _402611_402611 ; 
   reg __402611_402611;
   reg _402612_402612 ; 
   reg __402612_402612;
   reg _402613_402613 ; 
   reg __402613_402613;
   reg _402614_402614 ; 
   reg __402614_402614;
   reg _402615_402615 ; 
   reg __402615_402615;
   reg _402616_402616 ; 
   reg __402616_402616;
   reg _402617_402617 ; 
   reg __402617_402617;
   reg _402618_402618 ; 
   reg __402618_402618;
   reg _402619_402619 ; 
   reg __402619_402619;
   reg _402620_402620 ; 
   reg __402620_402620;
   reg _402621_402621 ; 
   reg __402621_402621;
   reg _402622_402622 ; 
   reg __402622_402622;
   reg _402623_402623 ; 
   reg __402623_402623;
   reg _402624_402624 ; 
   reg __402624_402624;
   reg _402625_402625 ; 
   reg __402625_402625;
   reg _402626_402626 ; 
   reg __402626_402626;
   reg _402627_402627 ; 
   reg __402627_402627;
   reg _402628_402628 ; 
   reg __402628_402628;
   reg _402629_402629 ; 
   reg __402629_402629;
   reg _402630_402630 ; 
   reg __402630_402630;
   reg _402631_402631 ; 
   reg __402631_402631;
   reg _402632_402632 ; 
   reg __402632_402632;
   reg _402633_402633 ; 
   reg __402633_402633;
   reg _402634_402634 ; 
   reg __402634_402634;
   reg _402635_402635 ; 
   reg __402635_402635;
   reg _402636_402636 ; 
   reg __402636_402636;
   reg _402637_402637 ; 
   reg __402637_402637;
   reg _402638_402638 ; 
   reg __402638_402638;
   reg _402639_402639 ; 
   reg __402639_402639;
   reg _402640_402640 ; 
   reg __402640_402640;
   reg _402641_402641 ; 
   reg __402641_402641;
   reg _402642_402642 ; 
   reg __402642_402642;
   reg _402643_402643 ; 
   reg __402643_402643;
   reg _402644_402644 ; 
   reg __402644_402644;
   reg _402645_402645 ; 
   reg __402645_402645;
   reg _402646_402646 ; 
   reg __402646_402646;
   reg _402647_402647 ; 
   reg __402647_402647;
   reg _402648_402648 ; 
   reg __402648_402648;
   reg _402649_402649 ; 
   reg __402649_402649;
   reg _402650_402650 ; 
   reg __402650_402650;
   reg _402651_402651 ; 
   reg __402651_402651;
   reg _402652_402652 ; 
   reg __402652_402652;
   reg _402653_402653 ; 
   reg __402653_402653;
   reg _402654_402654 ; 
   reg __402654_402654;
   reg _402655_402655 ; 
   reg __402655_402655;
   reg _402656_402656 ; 
   reg __402656_402656;
   reg _402657_402657 ; 
   reg __402657_402657;
   reg _402658_402658 ; 
   reg __402658_402658;
   reg _402659_402659 ; 
   reg __402659_402659;
   reg _402660_402660 ; 
   reg __402660_402660;
   reg _402661_402661 ; 
   reg __402661_402661;
   reg _402662_402662 ; 
   reg __402662_402662;
   reg _402663_402663 ; 
   reg __402663_402663;
   reg _402664_402664 ; 
   reg __402664_402664;
   reg _402665_402665 ; 
   reg __402665_402665;
   reg _402666_402666 ; 
   reg __402666_402666;
   reg _402667_402667 ; 
   reg __402667_402667;
   reg _402668_402668 ; 
   reg __402668_402668;
   reg _402669_402669 ; 
   reg __402669_402669;
   reg _402670_402670 ; 
   reg __402670_402670;
   reg _402671_402671 ; 
   reg __402671_402671;
   reg _402672_402672 ; 
   reg __402672_402672;
   reg _402673_402673 ; 
   reg __402673_402673;
   reg _402674_402674 ; 
   reg __402674_402674;
   reg _402675_402675 ; 
   reg __402675_402675;
   reg _402676_402676 ; 
   reg __402676_402676;
   reg _402677_402677 ; 
   reg __402677_402677;
   reg _402678_402678 ; 
   reg __402678_402678;
   reg _402679_402679 ; 
   reg __402679_402679;
   reg _402680_402680 ; 
   reg __402680_402680;
   reg _402681_402681 ; 
   reg __402681_402681;
   reg _402682_402682 ; 
   reg __402682_402682;
   reg _402683_402683 ; 
   reg __402683_402683;
   reg _402684_402684 ; 
   reg __402684_402684;
   reg _402685_402685 ; 
   reg __402685_402685;
   reg _402686_402686 ; 
   reg __402686_402686;
   reg _402687_402687 ; 
   reg __402687_402687;
   reg _402688_402688 ; 
   reg __402688_402688;
   reg _402689_402689 ; 
   reg __402689_402689;
   reg _402690_402690 ; 
   reg __402690_402690;
   reg _402691_402691 ; 
   reg __402691_402691;
   reg _402692_402692 ; 
   reg __402692_402692;
   reg _402693_402693 ; 
   reg __402693_402693;
   reg _402694_402694 ; 
   reg __402694_402694;
   reg _402695_402695 ; 
   reg __402695_402695;
   reg _402696_402696 ; 
   reg __402696_402696;
   reg _402697_402697 ; 
   reg __402697_402697;
   reg _402698_402698 ; 
   reg __402698_402698;
   reg _402699_402699 ; 
   reg __402699_402699;
   reg _402700_402700 ; 
   reg __402700_402700;
   reg _402701_402701 ; 
   reg __402701_402701;
   reg _402702_402702 ; 
   reg __402702_402702;
   reg _402703_402703 ; 
   reg __402703_402703;
   reg _402704_402704 ; 
   reg __402704_402704;
   reg _402705_402705 ; 
   reg __402705_402705;
   reg _402706_402706 ; 
   reg __402706_402706;
   reg _402707_402707 ; 
   reg __402707_402707;
   reg _402708_402708 ; 
   reg __402708_402708;
   reg _402709_402709 ; 
   reg __402709_402709;
   reg _402710_402710 ; 
   reg __402710_402710;
   reg _402711_402711 ; 
   reg __402711_402711;
   reg _402712_402712 ; 
   reg __402712_402712;
   reg _402713_402713 ; 
   reg __402713_402713;
   reg _402714_402714 ; 
   reg __402714_402714;
   reg _402715_402715 ; 
   reg __402715_402715;
   reg _402716_402716 ; 
   reg __402716_402716;
   reg _402717_402717 ; 
   reg __402717_402717;
   reg _402718_402718 ; 
   reg __402718_402718;
   reg _402719_402719 ; 
   reg __402719_402719;
   reg _402720_402720 ; 
   reg __402720_402720;
   reg _402721_402721 ; 
   reg __402721_402721;
   reg _402722_402722 ; 
   reg __402722_402722;
   reg _402723_402723 ; 
   reg __402723_402723;
   reg _402724_402724 ; 
   reg __402724_402724;
   reg _402725_402725 ; 
   reg __402725_402725;
   reg _402726_402726 ; 
   reg __402726_402726;
   reg _402727_402727 ; 
   reg __402727_402727;
   reg _402728_402728 ; 
   reg __402728_402728;
   reg _402729_402729 ; 
   reg __402729_402729;
   reg _402730_402730 ; 
   reg __402730_402730;
   reg _402731_402731 ; 
   reg __402731_402731;
   reg _402732_402732 ; 
   reg __402732_402732;
   reg _402733_402733 ; 
   reg __402733_402733;
   reg _402734_402734 ; 
   reg __402734_402734;
   reg _402735_402735 ; 
   reg __402735_402735;
   reg _402736_402736 ; 
   reg __402736_402736;
   reg _402737_402737 ; 
   reg __402737_402737;
   reg _402738_402738 ; 
   reg __402738_402738;
   reg _402739_402739 ; 
   reg __402739_402739;
   reg _402740_402740 ; 
   reg __402740_402740;
   reg _402741_402741 ; 
   reg __402741_402741;
   reg _402742_402742 ; 
   reg __402742_402742;
   reg _402743_402743 ; 
   reg __402743_402743;
   reg _402744_402744 ; 
   reg __402744_402744;
   reg _402745_402745 ; 
   reg __402745_402745;
   reg _402746_402746 ; 
   reg __402746_402746;
   reg _402747_402747 ; 
   reg __402747_402747;
   reg _402748_402748 ; 
   reg __402748_402748;
   reg _402749_402749 ; 
   reg __402749_402749;
   reg _402750_402750 ; 
   reg __402750_402750;
   reg _402751_402751 ; 
   reg __402751_402751;
   reg _402752_402752 ; 
   reg __402752_402752;
   reg _402753_402753 ; 
   reg __402753_402753;
   reg _402754_402754 ; 
   reg __402754_402754;
   reg _402755_402755 ; 
   reg __402755_402755;
   reg _402756_402756 ; 
   reg __402756_402756;
   reg _402757_402757 ; 
   reg __402757_402757;
   reg _402758_402758 ; 
   reg __402758_402758;
   reg _402759_402759 ; 
   reg __402759_402759;
   reg _402760_402760 ; 
   reg __402760_402760;
   reg _402761_402761 ; 
   reg __402761_402761;
   reg _402762_402762 ; 
   reg __402762_402762;
   reg _402763_402763 ; 
   reg __402763_402763;
   reg _402764_402764 ; 
   reg __402764_402764;
   reg _402765_402765 ; 
   reg __402765_402765;
   reg _402766_402766 ; 
   reg __402766_402766;
   reg _402767_402767 ; 
   reg __402767_402767;
   reg _402768_402768 ; 
   reg __402768_402768;
   reg _402769_402769 ; 
   reg __402769_402769;
   reg _402770_402770 ; 
   reg __402770_402770;
   reg _402771_402771 ; 
   reg __402771_402771;
   reg _402772_402772 ; 
   reg __402772_402772;
   reg _402773_402773 ; 
   reg __402773_402773;
   reg _402774_402774 ; 
   reg __402774_402774;
   reg _402775_402775 ; 
   reg __402775_402775;
   reg _402776_402776 ; 
   reg __402776_402776;
   reg _402777_402777 ; 
   reg __402777_402777;
   reg _402778_402778 ; 
   reg __402778_402778;
   reg _402779_402779 ; 
   reg __402779_402779;
   reg _402780_402780 ; 
   reg __402780_402780;
   reg _402781_402781 ; 
   reg __402781_402781;
   reg _402782_402782 ; 
   reg __402782_402782;
   reg _402783_402783 ; 
   reg __402783_402783;
   reg _402784_402784 ; 
   reg __402784_402784;
   reg _402785_402785 ; 
   reg __402785_402785;
   reg _402786_402786 ; 
   reg __402786_402786;
   reg _402787_402787 ; 
   reg __402787_402787;
   reg _402788_402788 ; 
   reg __402788_402788;
   reg _402789_402789 ; 
   reg __402789_402789;
   reg _402790_402790 ; 
   reg __402790_402790;
   reg _402791_402791 ; 
   reg __402791_402791;
   reg _402792_402792 ; 
   reg __402792_402792;
   reg _402793_402793 ; 
   reg __402793_402793;
   reg _402794_402794 ; 
   reg __402794_402794;
   reg _402795_402795 ; 
   reg __402795_402795;
   reg _402796_402796 ; 
   reg __402796_402796;
   reg _402797_402797 ; 
   reg __402797_402797;
   reg _402798_402798 ; 
   reg __402798_402798;
   reg _402799_402799 ; 
   reg __402799_402799;
   reg _402800_402800 ; 
   reg __402800_402800;
   reg _402801_402801 ; 
   reg __402801_402801;
   reg _402802_402802 ; 
   reg __402802_402802;
   reg _402803_402803 ; 
   reg __402803_402803;
   reg _402804_402804 ; 
   reg __402804_402804;
   reg _402805_402805 ; 
   reg __402805_402805;
   reg _402806_402806 ; 
   reg __402806_402806;
   reg _402807_402807 ; 
   reg __402807_402807;
   reg _402808_402808 ; 
   reg __402808_402808;
   reg _402809_402809 ; 
   reg __402809_402809;
   reg _402810_402810 ; 
   reg __402810_402810;
   reg _402811_402811 ; 
   reg __402811_402811;
   reg _402812_402812 ; 
   reg __402812_402812;
   reg _402813_402813 ; 
   reg __402813_402813;
   reg _402814_402814 ; 
   reg __402814_402814;
   reg _402815_402815 ; 
   reg __402815_402815;
   reg _402816_402816 ; 
   reg __402816_402816;
   reg _402817_402817 ; 
   reg __402817_402817;
   reg _402818_402818 ; 
   reg __402818_402818;
   reg _402819_402819 ; 
   reg __402819_402819;
   reg _402820_402820 ; 
   reg __402820_402820;
   reg _402821_402821 ; 
   reg __402821_402821;
   reg _402822_402822 ; 
   reg __402822_402822;
   reg _402823_402823 ; 
   reg __402823_402823;
   reg _402824_402824 ; 
   reg __402824_402824;
   reg _402825_402825 ; 
   reg __402825_402825;
   reg _402826_402826 ; 
   reg __402826_402826;
   reg _402827_402827 ; 
   reg __402827_402827;
   reg _402828_402828 ; 
   reg __402828_402828;
   reg _402829_402829 ; 
   reg __402829_402829;
   reg _402830_402830 ; 
   reg __402830_402830;
   reg _402831_402831 ; 
   reg __402831_402831;
   reg _402832_402832 ; 
   reg __402832_402832;
   reg _402833_402833 ; 
   reg __402833_402833;
   reg _402834_402834 ; 
   reg __402834_402834;
   reg _402835_402835 ; 
   reg __402835_402835;
   reg _402836_402836 ; 
   reg __402836_402836;
   reg _402837_402837 ; 
   reg __402837_402837;
   reg _402838_402838 ; 
   reg __402838_402838;
   reg _402839_402839 ; 
   reg __402839_402839;
   reg _402840_402840 ; 
   reg __402840_402840;
   reg _402841_402841 ; 
   reg __402841_402841;
   reg _402842_402842 ; 
   reg __402842_402842;
   reg _402843_402843 ; 
   reg __402843_402843;
   reg _402844_402844 ; 
   reg __402844_402844;
   reg _402845_402845 ; 
   reg __402845_402845;
   reg _402846_402846 ; 
   reg __402846_402846;
   reg _402847_402847 ; 
   reg __402847_402847;
   reg _402848_402848 ; 
   reg __402848_402848;
   reg _402849_402849 ; 
   reg __402849_402849;
   reg _402850_402850 ; 
   reg __402850_402850;
   reg _402851_402851 ; 
   reg __402851_402851;
   reg _402852_402852 ; 
   reg __402852_402852;
   reg _402853_402853 ; 
   reg __402853_402853;
   reg _402854_402854 ; 
   reg __402854_402854;
   reg _402855_402855 ; 
   reg __402855_402855;
   reg _402856_402856 ; 
   reg __402856_402856;
   reg _402857_402857 ; 
   reg __402857_402857;
   reg _402858_402858 ; 
   reg __402858_402858;
   reg _402859_402859 ; 
   reg __402859_402859;
   reg _402860_402860 ; 
   reg __402860_402860;
   reg _402861_402861 ; 
   reg __402861_402861;
   reg _402862_402862 ; 
   reg __402862_402862;
   reg _402863_402863 ; 
   reg __402863_402863;
   reg _402864_402864 ; 
   reg __402864_402864;
   reg _402865_402865 ; 
   reg __402865_402865;
   reg _402866_402866 ; 
   reg __402866_402866;
   reg _402867_402867 ; 
   reg __402867_402867;
   reg _402868_402868 ; 
   reg __402868_402868;
   reg _402869_402869 ; 
   reg __402869_402869;
   reg _402870_402870 ; 
   reg __402870_402870;
   reg _402871_402871 ; 
   reg __402871_402871;
   reg _402872_402872 ; 
   reg __402872_402872;
   reg _402873_402873 ; 
   reg __402873_402873;
   reg _402874_402874 ; 
   reg __402874_402874;
   reg _402875_402875 ; 
   reg __402875_402875;
   reg _402876_402876 ; 
   reg __402876_402876;
   reg _402877_402877 ; 
   reg __402877_402877;
   reg _402878_402878 ; 
   reg __402878_402878;
   reg _402879_402879 ; 
   reg __402879_402879;
   reg _402880_402880 ; 
   reg __402880_402880;
   reg _402881_402881 ; 
   reg __402881_402881;
   reg _402882_402882 ; 
   reg __402882_402882;
   reg _402883_402883 ; 
   reg __402883_402883;
   reg _402884_402884 ; 
   reg __402884_402884;
   reg _402885_402885 ; 
   reg __402885_402885;
   reg _402886_402886 ; 
   reg __402886_402886;
   reg _402887_402887 ; 
   reg __402887_402887;
   reg _402888_402888 ; 
   reg __402888_402888;
   reg _402889_402889 ; 
   reg __402889_402889;
   reg _402890_402890 ; 
   reg __402890_402890;
   reg _402891_402891 ; 
   reg __402891_402891;
   reg _402892_402892 ; 
   reg __402892_402892;
   reg _402893_402893 ; 
   reg __402893_402893;
   reg _402894_402894 ; 
   reg __402894_402894;
   reg _402895_402895 ; 
   reg __402895_402895;
   reg _402896_402896 ; 
   reg __402896_402896;
   reg _402897_402897 ; 
   reg __402897_402897;
   reg _402898_402898 ; 
   reg __402898_402898;
   reg _402899_402899 ; 
   reg __402899_402899;
   reg _402900_402900 ; 
   reg __402900_402900;
   reg _402901_402901 ; 
   reg __402901_402901;
   reg _402902_402902 ; 
   reg __402902_402902;
   reg _402903_402903 ; 
   reg __402903_402903;
   reg _402904_402904 ; 
   reg __402904_402904;
   reg _402905_402905 ; 
   reg __402905_402905;
   reg _402906_402906 ; 
   reg __402906_402906;
   reg _402907_402907 ; 
   reg __402907_402907;
   reg _402908_402908 ; 
   reg __402908_402908;
   reg _402909_402909 ; 
   reg __402909_402909;
   reg _402910_402910 ; 
   reg __402910_402910;
   reg _402911_402911 ; 
   reg __402911_402911;
   reg _402912_402912 ; 
   reg __402912_402912;
   reg _402913_402913 ; 
   reg __402913_402913;
   reg _402914_402914 ; 
   reg __402914_402914;
   reg _402915_402915 ; 
   reg __402915_402915;
   reg _402916_402916 ; 
   reg __402916_402916;
   reg _402917_402917 ; 
   reg __402917_402917;
   reg _402918_402918 ; 
   reg __402918_402918;
   reg _402919_402919 ; 
   reg __402919_402919;
   reg _402920_402920 ; 
   reg __402920_402920;
   reg _402921_402921 ; 
   reg __402921_402921;
   reg _402922_402922 ; 
   reg __402922_402922;
   reg _402923_402923 ; 
   reg __402923_402923;
   reg _402924_402924 ; 
   reg __402924_402924;
   reg _402925_402925 ; 
   reg __402925_402925;
   reg _402926_402926 ; 
   reg __402926_402926;
   reg _402927_402927 ; 
   reg __402927_402927;
   reg _402928_402928 ; 
   reg __402928_402928;
   reg _402929_402929 ; 
   reg __402929_402929;
   reg _402930_402930 ; 
   reg __402930_402930;
   reg _402931_402931 ; 
   reg __402931_402931;
   reg _402932_402932 ; 
   reg __402932_402932;
   reg _402933_402933 ; 
   reg __402933_402933;
   reg _402934_402934 ; 
   reg __402934_402934;
   reg _402935_402935 ; 
   reg __402935_402935;
   reg _402936_402936 ; 
   reg __402936_402936;
   reg _402937_402937 ; 
   reg __402937_402937;
   reg _402938_402938 ; 
   reg __402938_402938;
   reg _402939_402939 ; 
   reg __402939_402939;
   reg _402940_402940 ; 
   reg __402940_402940;
   reg _402941_402941 ; 
   reg __402941_402941;
   reg _402942_402942 ; 
   reg __402942_402942;
   reg _402943_402943 ; 
   reg __402943_402943;
   reg _402944_402944 ; 
   reg __402944_402944;
   reg _402945_402945 ; 
   reg __402945_402945;
   reg _402946_402946 ; 
   reg __402946_402946;
   reg _402947_402947 ; 
   reg __402947_402947;
   reg _402948_402948 ; 
   reg __402948_402948;
   reg _402949_402949 ; 
   reg __402949_402949;
   reg _402950_402950 ; 
   reg __402950_402950;
   reg _402951_402951 ; 
   reg __402951_402951;
   reg _402952_402952 ; 
   reg __402952_402952;
   reg _402953_402953 ; 
   reg __402953_402953;
   reg _402954_402954 ; 
   reg __402954_402954;
   reg _402955_402955 ; 
   reg __402955_402955;
   reg _402956_402956 ; 
   reg __402956_402956;
   reg _402957_402957 ; 
   reg __402957_402957;
   reg _402958_402958 ; 
   reg __402958_402958;
   reg _402959_402959 ; 
   reg __402959_402959;
   reg _402960_402960 ; 
   reg __402960_402960;
   reg _402961_402961 ; 
   reg __402961_402961;
   reg _402962_402962 ; 
   reg __402962_402962;
   reg _402963_402963 ; 
   reg __402963_402963;
   reg _402964_402964 ; 
   reg __402964_402964;
   reg _402965_402965 ; 
   reg __402965_402965;
   reg _402966_402966 ; 
   reg __402966_402966;
   reg _402967_402967 ; 
   reg __402967_402967;
   reg _402968_402968 ; 
   reg __402968_402968;
   reg _402969_402969 ; 
   reg __402969_402969;
   reg _402970_402970 ; 
   reg __402970_402970;
   reg _402971_402971 ; 
   reg __402971_402971;
   reg _402972_402972 ; 
   reg __402972_402972;
   reg _402973_402973 ; 
   reg __402973_402973;
   reg _402974_402974 ; 
   reg __402974_402974;
   reg _402975_402975 ; 
   reg __402975_402975;
   reg _402976_402976 ; 
   reg __402976_402976;
   reg _402977_402977 ; 
   reg __402977_402977;
   reg _402978_402978 ; 
   reg __402978_402978;
   reg _402979_402979 ; 
   reg __402979_402979;
   reg _402980_402980 ; 
   reg __402980_402980;
   reg _402981_402981 ; 
   reg __402981_402981;
   reg _402982_402982 ; 
   reg __402982_402982;
   reg _402983_402983 ; 
   reg __402983_402983;
   reg _402984_402984 ; 
   reg __402984_402984;
   reg _402985_402985 ; 
   reg __402985_402985;
   reg _402986_402986 ; 
   reg __402986_402986;
   reg _402987_402987 ; 
   reg __402987_402987;
   reg _402988_402988 ; 
   reg __402988_402988;
   reg _402989_402989 ; 
   reg __402989_402989;
   reg _402990_402990 ; 
   reg __402990_402990;
   reg _402991_402991 ; 
   reg __402991_402991;
   reg _402992_402992 ; 
   reg __402992_402992;
   reg _402993_402993 ; 
   reg __402993_402993;
   reg _402994_402994 ; 
   reg __402994_402994;
   reg _402995_402995 ; 
   reg __402995_402995;
   reg _402996_402996 ; 
   reg __402996_402996;
   reg _402997_402997 ; 
   reg __402997_402997;
   reg _402998_402998 ; 
   reg __402998_402998;
   reg _402999_402999 ; 
   reg __402999_402999;
   reg _403000_403000 ; 
   reg __403000_403000;
   reg _403001_403001 ; 
   reg __403001_403001;
   reg _403002_403002 ; 
   reg __403002_403002;
   reg _403003_403003 ; 
   reg __403003_403003;
   reg _403004_403004 ; 
   reg __403004_403004;
   reg _403005_403005 ; 
   reg __403005_403005;
   reg _403006_403006 ; 
   reg __403006_403006;
   reg _403007_403007 ; 
   reg __403007_403007;
   reg _403008_403008 ; 
   reg __403008_403008;
   reg _403009_403009 ; 
   reg __403009_403009;
   reg _403010_403010 ; 
   reg __403010_403010;
   reg _403011_403011 ; 
   reg __403011_403011;
   reg _403012_403012 ; 
   reg __403012_403012;
   reg _403013_403013 ; 
   reg __403013_403013;
   reg _403014_403014 ; 
   reg __403014_403014;
   reg _403015_403015 ; 
   reg __403015_403015;
   reg _403016_403016 ; 
   reg __403016_403016;
   reg _403017_403017 ; 
   reg __403017_403017;
   reg _403018_403018 ; 
   reg __403018_403018;
   reg _403019_403019 ; 
   reg __403019_403019;
   reg _403020_403020 ; 
   reg __403020_403020;
   reg _403021_403021 ; 
   reg __403021_403021;
   reg _403022_403022 ; 
   reg __403022_403022;
   reg _403023_403023 ; 
   reg __403023_403023;
   reg _403024_403024 ; 
   reg __403024_403024;
   reg _403025_403025 ; 
   reg __403025_403025;
   reg _403026_403026 ; 
   reg __403026_403026;
   reg _403027_403027 ; 
   reg __403027_403027;
   reg _403028_403028 ; 
   reg __403028_403028;
   reg _403029_403029 ; 
   reg __403029_403029;
   reg _403030_403030 ; 
   reg __403030_403030;
   reg _403031_403031 ; 
   reg __403031_403031;
   reg _403032_403032 ; 
   reg __403032_403032;
   reg _403033_403033 ; 
   reg __403033_403033;
   reg _403034_403034 ; 
   reg __403034_403034;
   reg _403035_403035 ; 
   reg __403035_403035;
   reg _403036_403036 ; 
   reg __403036_403036;
   reg _403037_403037 ; 
   reg __403037_403037;
   reg _403038_403038 ; 
   reg __403038_403038;
   reg _403039_403039 ; 
   reg __403039_403039;
   reg _403040_403040 ; 
   reg __403040_403040;
   reg _403041_403041 ; 
   reg __403041_403041;
   reg _403042_403042 ; 
   reg __403042_403042;
   reg _403043_403043 ; 
   reg __403043_403043;
   reg _403044_403044 ; 
   reg __403044_403044;
   reg _403045_403045 ; 
   reg __403045_403045;
   reg _403046_403046 ; 
   reg __403046_403046;
   reg _403047_403047 ; 
   reg __403047_403047;
   reg _403048_403048 ; 
   reg __403048_403048;
   reg _403049_403049 ; 
   reg __403049_403049;
   reg _403050_403050 ; 
   reg __403050_403050;
   reg _403051_403051 ; 
   reg __403051_403051;
   reg _403052_403052 ; 
   reg __403052_403052;
   reg _403053_403053 ; 
   reg __403053_403053;
   reg _403054_403054 ; 
   reg __403054_403054;
   reg _403055_403055 ; 
   reg __403055_403055;
   reg _403056_403056 ; 
   reg __403056_403056;
   reg _403057_403057 ; 
   reg __403057_403057;
   reg _403058_403058 ; 
   reg __403058_403058;
   reg _403059_403059 ; 
   reg __403059_403059;
   reg _403060_403060 ; 
   reg __403060_403060;
   reg _403061_403061 ; 
   reg __403061_403061;
   reg _403062_403062 ; 
   reg __403062_403062;
   reg _403063_403063 ; 
   reg __403063_403063;
   reg _403064_403064 ; 
   reg __403064_403064;
   reg _403065_403065 ; 
   reg __403065_403065;
   reg _403066_403066 ; 
   reg __403066_403066;
   reg _403067_403067 ; 
   reg __403067_403067;
   reg _403068_403068 ; 
   reg __403068_403068;
   reg _403069_403069 ; 
   reg __403069_403069;
   reg _403070_403070 ; 
   reg __403070_403070;
   reg _403071_403071 ; 
   reg __403071_403071;
   reg _403072_403072 ; 
   reg __403072_403072;
   reg _403073_403073 ; 
   reg __403073_403073;
   reg _403074_403074 ; 
   reg __403074_403074;
   reg _403075_403075 ; 
   reg __403075_403075;
   reg _403076_403076 ; 
   reg __403076_403076;
   reg _403077_403077 ; 
   reg __403077_403077;
   reg _403078_403078 ; 
   reg __403078_403078;
   reg _403079_403079 ; 
   reg __403079_403079;
   reg _403080_403080 ; 
   reg __403080_403080;
   reg _403081_403081 ; 
   reg __403081_403081;
   reg _403082_403082 ; 
   reg __403082_403082;
   reg _403083_403083 ; 
   reg __403083_403083;
   reg _403084_403084 ; 
   reg __403084_403084;
   reg _403085_403085 ; 
   reg __403085_403085;
   reg _403086_403086 ; 
   reg __403086_403086;
   reg _403087_403087 ; 
   reg __403087_403087;
   reg _403088_403088 ; 
   reg __403088_403088;
   reg _403089_403089 ; 
   reg __403089_403089;
   reg _403090_403090 ; 
   reg __403090_403090;
   reg _403091_403091 ; 
   reg __403091_403091;
   reg _403092_403092 ; 
   reg __403092_403092;
   reg _403093_403093 ; 
   reg __403093_403093;
   reg _403094_403094 ; 
   reg __403094_403094;
   reg _403095_403095 ; 
   reg __403095_403095;
   reg _403096_403096 ; 
   reg __403096_403096;
   reg _403097_403097 ; 
   reg __403097_403097;
   reg _403098_403098 ; 
   reg __403098_403098;
   reg _403099_403099 ; 
   reg __403099_403099;
   reg _403100_403100 ; 
   reg __403100_403100;
   reg _403101_403101 ; 
   reg __403101_403101;
   reg _403102_403102 ; 
   reg __403102_403102;
   reg _403103_403103 ; 
   reg __403103_403103;
   reg _403104_403104 ; 
   reg __403104_403104;
   reg _403105_403105 ; 
   reg __403105_403105;
   reg _403106_403106 ; 
   reg __403106_403106;
   reg _403107_403107 ; 
   reg __403107_403107;
   reg _403108_403108 ; 
   reg __403108_403108;
   reg _403109_403109 ; 
   reg __403109_403109;
   reg _403110_403110 ; 
   reg __403110_403110;
   reg _403111_403111 ; 
   reg __403111_403111;
   reg _403112_403112 ; 
   reg __403112_403112;
   reg _403113_403113 ; 
   reg __403113_403113;
   reg _403114_403114 ; 
   reg __403114_403114;
   reg _403115_403115 ; 
   reg __403115_403115;
   reg _403116_403116 ; 
   reg __403116_403116;
   reg _403117_403117 ; 
   reg __403117_403117;
   reg _403118_403118 ; 
   reg __403118_403118;
   reg _403119_403119 ; 
   reg __403119_403119;
   reg _403120_403120 ; 
   reg __403120_403120;
   reg _403121_403121 ; 
   reg __403121_403121;
   reg _403122_403122 ; 
   reg __403122_403122;
   reg _403123_403123 ; 
   reg __403123_403123;
   reg _403124_403124 ; 
   reg __403124_403124;
   reg _403125_403125 ; 
   reg __403125_403125;
   reg _403126_403126 ; 
   reg __403126_403126;
   reg _403127_403127 ; 
   reg __403127_403127;
   reg _403128_403128 ; 
   reg __403128_403128;
   reg _403129_403129 ; 
   reg __403129_403129;
   reg _403130_403130 ; 
   reg __403130_403130;
   reg _403131_403131 ; 
   reg __403131_403131;
   reg _403132_403132 ; 
   reg __403132_403132;
   reg _403133_403133 ; 
   reg __403133_403133;
   reg _403134_403134 ; 
   reg __403134_403134;
   reg _403135_403135 ; 
   reg __403135_403135;
   reg _403136_403136 ; 
   reg __403136_403136;
   reg _403137_403137 ; 
   reg __403137_403137;
   reg _403138_403138 ; 
   reg __403138_403138;
   reg _403139_403139 ; 
   reg __403139_403139;
   reg _403140_403140 ; 
   reg __403140_403140;
   reg _403141_403141 ; 
   reg __403141_403141;
   reg _403142_403142 ; 
   reg __403142_403142;
   reg _403143_403143 ; 
   reg __403143_403143;
   reg _403144_403144 ; 
   reg __403144_403144;
   reg _403145_403145 ; 
   reg __403145_403145;
   reg _403146_403146 ; 
   reg __403146_403146;
   reg _403147_403147 ; 
   reg __403147_403147;
   reg _403148_403148 ; 
   reg __403148_403148;
   reg _403149_403149 ; 
   reg __403149_403149;
   reg _403150_403150 ; 
   reg __403150_403150;
   reg _403151_403151 ; 
   reg __403151_403151;
   reg _403152_403152 ; 
   reg __403152_403152;
   reg _403153_403153 ; 
   reg __403153_403153;
   reg _403154_403154 ; 
   reg __403154_403154;
   reg _403155_403155 ; 
   reg __403155_403155;
   reg _403156_403156 ; 
   reg __403156_403156;
   reg _403157_403157 ; 
   reg __403157_403157;
   reg _403158_403158 ; 
   reg __403158_403158;
   reg _403159_403159 ; 
   reg __403159_403159;
   reg _403160_403160 ; 
   reg __403160_403160;
   reg _403161_403161 ; 
   reg __403161_403161;
   reg _403162_403162 ; 
   reg __403162_403162;
   reg _403163_403163 ; 
   reg __403163_403163;
   reg _403164_403164 ; 
   reg __403164_403164;
   reg _403165_403165 ; 
   reg __403165_403165;
   reg _403166_403166 ; 
   reg __403166_403166;
   reg _403167_403167 ; 
   reg __403167_403167;
   reg _403168_403168 ; 
   reg __403168_403168;
   reg _403169_403169 ; 
   reg __403169_403169;
   reg _403170_403170 ; 
   reg __403170_403170;
   reg _403171_403171 ; 
   reg __403171_403171;
   reg _403172_403172 ; 
   reg __403172_403172;
   reg _403173_403173 ; 
   reg __403173_403173;
   reg _403174_403174 ; 
   reg __403174_403174;
   reg _403175_403175 ; 
   reg __403175_403175;
   reg _403176_403176 ; 
   reg __403176_403176;
   reg _403177_403177 ; 
   reg __403177_403177;
   reg _403178_403178 ; 
   reg __403178_403178;
   reg _403179_403179 ; 
   reg __403179_403179;
   reg _403180_403180 ; 
   reg __403180_403180;
   reg _403181_403181 ; 
   reg __403181_403181;
   reg _403182_403182 ; 
   reg __403182_403182;
   reg _403183_403183 ; 
   reg __403183_403183;
   reg _403184_403184 ; 
   reg __403184_403184;
   reg _403185_403185 ; 
   reg __403185_403185;
   reg _403186_403186 ; 
   reg __403186_403186;
   reg _403187_403187 ; 
   reg __403187_403187;
   reg _403188_403188 ; 
   reg __403188_403188;
   reg _403189_403189 ; 
   reg __403189_403189;
   reg _403190_403190 ; 
   reg __403190_403190;
   reg _403191_403191 ; 
   reg __403191_403191;
   reg _403192_403192 ; 
   reg __403192_403192;
   reg _403193_403193 ; 
   reg __403193_403193;
   reg _403194_403194 ; 
   reg __403194_403194;
   reg _403195_403195 ; 
   reg __403195_403195;
   reg _403196_403196 ; 
   reg __403196_403196;
   reg _403197_403197 ; 
   reg __403197_403197;
   reg _403198_403198 ; 
   reg __403198_403198;
   reg _403199_403199 ; 
   reg __403199_403199;
   reg _403200_403200 ; 
   reg __403200_403200;
   reg _403201_403201 ; 
   reg __403201_403201;
   reg _403202_403202 ; 
   reg __403202_403202;
   reg _403203_403203 ; 
   reg __403203_403203;
   reg _403204_403204 ; 
   reg __403204_403204;
   reg _403205_403205 ; 
   reg __403205_403205;
   reg _403206_403206 ; 
   reg __403206_403206;
   reg _403207_403207 ; 
   reg __403207_403207;
   reg _403208_403208 ; 
   reg __403208_403208;
   reg _403209_403209 ; 
   reg __403209_403209;
   reg _403210_403210 ; 
   reg __403210_403210;
   reg _403211_403211 ; 
   reg __403211_403211;
   reg _403212_403212 ; 
   reg __403212_403212;
   reg _403213_403213 ; 
   reg __403213_403213;
   reg _403214_403214 ; 
   reg __403214_403214;
   reg _403215_403215 ; 
   reg __403215_403215;
   reg _403216_403216 ; 
   reg __403216_403216;
   reg _403217_403217 ; 
   reg __403217_403217;
   reg _403218_403218 ; 
   reg __403218_403218;
   reg _403219_403219 ; 
   reg __403219_403219;
   reg _403220_403220 ; 
   reg __403220_403220;
   reg _403221_403221 ; 
   reg __403221_403221;
   reg _403222_403222 ; 
   reg __403222_403222;
   reg _403223_403223 ; 
   reg __403223_403223;
   reg _403224_403224 ; 
   reg __403224_403224;
   reg _403225_403225 ; 
   reg __403225_403225;
   reg _403226_403226 ; 
   reg __403226_403226;
   reg _403227_403227 ; 
   reg __403227_403227;
   reg _403228_403228 ; 
   reg __403228_403228;
   reg _403229_403229 ; 
   reg __403229_403229;
   reg _403230_403230 ; 
   reg __403230_403230;
   reg _403231_403231 ; 
   reg __403231_403231;
   reg _403232_403232 ; 
   reg __403232_403232;
   reg _403233_403233 ; 
   reg __403233_403233;
   reg _403234_403234 ; 
   reg __403234_403234;
   reg _403235_403235 ; 
   reg __403235_403235;
   reg _403236_403236 ; 
   reg __403236_403236;
   reg _403237_403237 ; 
   reg __403237_403237;
   reg _403238_403238 ; 
   reg __403238_403238;
   reg _403239_403239 ; 
   reg __403239_403239;
   reg _403240_403240 ; 
   reg __403240_403240;
   reg _403241_403241 ; 
   reg __403241_403241;
   reg _403242_403242 ; 
   reg __403242_403242;
   reg _403243_403243 ; 
   reg __403243_403243;
   reg _403244_403244 ; 
   reg __403244_403244;
   reg _403245_403245 ; 
   reg __403245_403245;
   reg _403246_403246 ; 
   reg __403246_403246;
   reg _403247_403247 ; 
   reg __403247_403247;
   reg _403248_403248 ; 
   reg __403248_403248;
   reg _403249_403249 ; 
   reg __403249_403249;
   reg _403250_403250 ; 
   reg __403250_403250;
   reg _403251_403251 ; 
   reg __403251_403251;
   reg _403252_403252 ; 
   reg __403252_403252;
   reg _403253_403253 ; 
   reg __403253_403253;
   reg _403254_403254 ; 
   reg __403254_403254;
   reg _403255_403255 ; 
   reg __403255_403255;
   reg _403256_403256 ; 
   reg __403256_403256;
   reg _403257_403257 ; 
   reg __403257_403257;
   reg _403258_403258 ; 
   reg __403258_403258;
   reg _403259_403259 ; 
   reg __403259_403259;
   reg _403260_403260 ; 
   reg __403260_403260;
   reg _403261_403261 ; 
   reg __403261_403261;
   reg _403262_403262 ; 
   reg __403262_403262;
   reg _403263_403263 ; 
   reg __403263_403263;
   reg _403264_403264 ; 
   reg __403264_403264;
   reg _403265_403265 ; 
   reg __403265_403265;
   reg _403266_403266 ; 
   reg __403266_403266;
   reg _403267_403267 ; 
   reg __403267_403267;
   reg _403268_403268 ; 
   reg __403268_403268;
   reg _403269_403269 ; 
   reg __403269_403269;
   reg _403270_403270 ; 
   reg __403270_403270;
   reg _403271_403271 ; 
   reg __403271_403271;
   reg _403272_403272 ; 
   reg __403272_403272;
   reg _403273_403273 ; 
   reg __403273_403273;
   reg _403274_403274 ; 
   reg __403274_403274;
   reg _403275_403275 ; 
   reg __403275_403275;
   reg _403276_403276 ; 
   reg __403276_403276;
   reg _403277_403277 ; 
   reg __403277_403277;
   reg _403278_403278 ; 
   reg __403278_403278;
   reg _403279_403279 ; 
   reg __403279_403279;
   reg _403280_403280 ; 
   reg __403280_403280;
   reg _403281_403281 ; 
   reg __403281_403281;
   reg _403282_403282 ; 
   reg __403282_403282;
   reg _403283_403283 ; 
   reg __403283_403283;
   reg _403284_403284 ; 
   reg __403284_403284;
   reg _403285_403285 ; 
   reg __403285_403285;
   reg _403286_403286 ; 
   reg __403286_403286;
   reg _403287_403287 ; 
   reg __403287_403287;
   reg _403288_403288 ; 
   reg __403288_403288;
   reg _403289_403289 ; 
   reg __403289_403289;
   reg _403290_403290 ; 
   reg __403290_403290;
   reg _403291_403291 ; 
   reg __403291_403291;
   reg _403292_403292 ; 
   reg __403292_403292;
   reg _403293_403293 ; 
   reg __403293_403293;
   reg _403294_403294 ; 
   reg __403294_403294;
   reg _403295_403295 ; 
   reg __403295_403295;
   reg _403296_403296 ; 
   reg __403296_403296;
   reg _403297_403297 ; 
   reg __403297_403297;
   reg _403298_403298 ; 
   reg __403298_403298;
   reg _403299_403299 ; 
   reg __403299_403299;
   reg _403300_403300 ; 
   reg __403300_403300;
   reg _403301_403301 ; 
   reg __403301_403301;
   reg _403302_403302 ; 
   reg __403302_403302;
   reg _403303_403303 ; 
   reg __403303_403303;
   reg _403304_403304 ; 
   reg __403304_403304;
   reg _403305_403305 ; 
   reg __403305_403305;
   reg _403306_403306 ; 
   reg __403306_403306;
   reg _403307_403307 ; 
   reg __403307_403307;
   reg _403308_403308 ; 
   reg __403308_403308;
   reg _403309_403309 ; 
   reg __403309_403309;
   reg _403310_403310 ; 
   reg __403310_403310;
   reg _403311_403311 ; 
   reg __403311_403311;
   reg _403312_403312 ; 
   reg __403312_403312;
   reg _403313_403313 ; 
   reg __403313_403313;
   reg _403314_403314 ; 
   reg __403314_403314;
   reg _403315_403315 ; 
   reg __403315_403315;
   reg _403316_403316 ; 
   reg __403316_403316;
   reg _403317_403317 ; 
   reg __403317_403317;
   reg _403318_403318 ; 
   reg __403318_403318;
   reg _403319_403319 ; 
   reg __403319_403319;
   reg _403320_403320 ; 
   reg __403320_403320;
   reg _403321_403321 ; 
   reg __403321_403321;
   reg _403322_403322 ; 
   reg __403322_403322;
   reg _403323_403323 ; 
   reg __403323_403323;
   reg _403324_403324 ; 
   reg __403324_403324;
   reg _403325_403325 ; 
   reg __403325_403325;
   reg _403326_403326 ; 
   reg __403326_403326;
   reg _403327_403327 ; 
   reg __403327_403327;
   reg _403328_403328 ; 
   reg __403328_403328;
   reg _403329_403329 ; 
   reg __403329_403329;
   reg _403330_403330 ; 
   reg __403330_403330;
   reg _403331_403331 ; 
   reg __403331_403331;
   reg _403332_403332 ; 
   reg __403332_403332;
   reg _403333_403333 ; 
   reg __403333_403333;
   reg _403334_403334 ; 
   reg __403334_403334;
   reg _403335_403335 ; 
   reg __403335_403335;
   reg _403336_403336 ; 
   reg __403336_403336;
   reg _403337_403337 ; 
   reg __403337_403337;
   reg _403338_403338 ; 
   reg __403338_403338;
   reg _403339_403339 ; 
   reg __403339_403339;
   reg _403340_403340 ; 
   reg __403340_403340;
   reg _403341_403341 ; 
   reg __403341_403341;
   reg _403342_403342 ; 
   reg __403342_403342;
   reg _403343_403343 ; 
   reg __403343_403343;
   reg _403344_403344 ; 
   reg __403344_403344;
   reg _403345_403345 ; 
   reg __403345_403345;
   reg _403346_403346 ; 
   reg __403346_403346;
   reg _403347_403347 ; 
   reg __403347_403347;
   reg _403348_403348 ; 
   reg __403348_403348;
   reg _403349_403349 ; 
   reg __403349_403349;
   reg _403350_403350 ; 
   reg __403350_403350;
   reg _403351_403351 ; 
   reg __403351_403351;
   reg _403352_403352 ; 
   reg __403352_403352;
   reg _403353_403353 ; 
   reg __403353_403353;
   reg _403354_403354 ; 
   reg __403354_403354;
   reg _403355_403355 ; 
   reg __403355_403355;
   reg _403356_403356 ; 
   reg __403356_403356;
   reg _403357_403357 ; 
   reg __403357_403357;
   reg _403358_403358 ; 
   reg __403358_403358;
   reg _403359_403359 ; 
   reg __403359_403359;
   reg _403360_403360 ; 
   reg __403360_403360;
   reg _403361_403361 ; 
   reg __403361_403361;
   reg _403362_403362 ; 
   reg __403362_403362;
   reg _403363_403363 ; 
   reg __403363_403363;
   reg _403364_403364 ; 
   reg __403364_403364;
   reg _403365_403365 ; 
   reg __403365_403365;
   reg _403366_403366 ; 
   reg __403366_403366;
   reg _403367_403367 ; 
   reg __403367_403367;
   reg _403368_403368 ; 
   reg __403368_403368;
   reg _403369_403369 ; 
   reg __403369_403369;
   reg _403370_403370 ; 
   reg __403370_403370;
   reg _403371_403371 ; 
   reg __403371_403371;
   reg _403372_403372 ; 
   reg __403372_403372;
   reg _403373_403373 ; 
   reg __403373_403373;
   reg _403374_403374 ; 
   reg __403374_403374;
   reg _403375_403375 ; 
   reg __403375_403375;
   reg _403376_403376 ; 
   reg __403376_403376;
   reg _403377_403377 ; 
   reg __403377_403377;
   reg _403378_403378 ; 
   reg __403378_403378;
   reg _403379_403379 ; 
   reg __403379_403379;
   reg _403380_403380 ; 
   reg __403380_403380;
   reg _403381_403381 ; 
   reg __403381_403381;
   reg _403382_403382 ; 
   reg __403382_403382;
   reg _403383_403383 ; 
   reg __403383_403383;
   reg _403384_403384 ; 
   reg __403384_403384;
   reg _403385_403385 ; 
   reg __403385_403385;
   reg _403386_403386 ; 
   reg __403386_403386;
   reg _403387_403387 ; 
   reg __403387_403387;
   reg _403388_403388 ; 
   reg __403388_403388;
   reg _403389_403389 ; 
   reg __403389_403389;
   reg _403390_403390 ; 
   reg __403390_403390;
   reg _403391_403391 ; 
   reg __403391_403391;
   reg _403392_403392 ; 
   reg __403392_403392;
   reg _403393_403393 ; 
   reg __403393_403393;
   reg _403394_403394 ; 
   reg __403394_403394;
   reg _403395_403395 ; 
   reg __403395_403395;
   reg _403396_403396 ; 
   reg __403396_403396;
   reg _403397_403397 ; 
   reg __403397_403397;
   reg _403398_403398 ; 
   reg __403398_403398;
   reg _403399_403399 ; 
   reg __403399_403399;
   reg _403400_403400 ; 
   reg __403400_403400;
   reg _403401_403401 ; 
   reg __403401_403401;
   reg _403402_403402 ; 
   reg __403402_403402;
   reg _403403_403403 ; 
   reg __403403_403403;
   reg _403404_403404 ; 
   reg __403404_403404;
   reg _403405_403405 ; 
   reg __403405_403405;
   reg _403406_403406 ; 
   reg __403406_403406;
   reg _403407_403407 ; 
   reg __403407_403407;
   reg _403408_403408 ; 
   reg __403408_403408;
   reg _403409_403409 ; 
   reg __403409_403409;
   reg _403410_403410 ; 
   reg __403410_403410;
   reg _403411_403411 ; 
   reg __403411_403411;
   reg _403412_403412 ; 
   reg __403412_403412;
   reg _403413_403413 ; 
   reg __403413_403413;
   reg _403414_403414 ; 
   reg __403414_403414;
   reg _403415_403415 ; 
   reg __403415_403415;
   reg _403416_403416 ; 
   reg __403416_403416;
   reg _403417_403417 ; 
   reg __403417_403417;
   reg _403418_403418 ; 
   reg __403418_403418;
   reg _403419_403419 ; 
   reg __403419_403419;
   reg _403420_403420 ; 
   reg __403420_403420;
   reg _403421_403421 ; 
   reg __403421_403421;
   reg _403422_403422 ; 
   reg __403422_403422;
   reg _403423_403423 ; 
   reg __403423_403423;
   reg _403424_403424 ; 
   reg __403424_403424;
   reg _403425_403425 ; 
   reg __403425_403425;
   reg _403426_403426 ; 
   reg __403426_403426;
   reg _403427_403427 ; 
   reg __403427_403427;
   reg _403428_403428 ; 
   reg __403428_403428;
   reg _403429_403429 ; 
   reg __403429_403429;
   reg _403430_403430 ; 
   reg __403430_403430;
   reg _403431_403431 ; 
   reg __403431_403431;
   reg _403432_403432 ; 
   reg __403432_403432;
   reg _403433_403433 ; 
   reg __403433_403433;
   reg _403434_403434 ; 
   reg __403434_403434;
   reg _403435_403435 ; 
   reg __403435_403435;
   reg _403436_403436 ; 
   reg __403436_403436;
   reg _403437_403437 ; 
   reg __403437_403437;
   reg _403438_403438 ; 
   reg __403438_403438;
   reg _403439_403439 ; 
   reg __403439_403439;
   reg _403440_403440 ; 
   reg __403440_403440;
   reg _403441_403441 ; 
   reg __403441_403441;
   reg _403442_403442 ; 
   reg __403442_403442;
   reg _403443_403443 ; 
   reg __403443_403443;
   reg _403444_403444 ; 
   reg __403444_403444;
   reg _403445_403445 ; 
   reg __403445_403445;
   reg _403446_403446 ; 
   reg __403446_403446;
   reg _403447_403447 ; 
   reg __403447_403447;
   reg _403448_403448 ; 
   reg __403448_403448;
   reg _403449_403449 ; 
   reg __403449_403449;
   reg _403450_403450 ; 
   reg __403450_403450;
   reg _403451_403451 ; 
   reg __403451_403451;
   reg _403452_403452 ; 
   reg __403452_403452;
   reg _403453_403453 ; 
   reg __403453_403453;
   reg _403454_403454 ; 
   reg __403454_403454;
   reg _403455_403455 ; 
   reg __403455_403455;
   reg _403456_403456 ; 
   reg __403456_403456;
   reg _403457_403457 ; 
   reg __403457_403457;
   reg _403458_403458 ; 
   reg __403458_403458;
   reg _403459_403459 ; 
   reg __403459_403459;
   reg _403460_403460 ; 
   reg __403460_403460;
   reg _403461_403461 ; 
   reg __403461_403461;
   reg _403462_403462 ; 
   reg __403462_403462;
   reg _403463_403463 ; 
   reg __403463_403463;
   reg _403464_403464 ; 
   reg __403464_403464;
   reg _403465_403465 ; 
   reg __403465_403465;
   reg _403466_403466 ; 
   reg __403466_403466;
   reg _403467_403467 ; 
   reg __403467_403467;
   reg _403468_403468 ; 
   reg __403468_403468;
   reg _403469_403469 ; 
   reg __403469_403469;
   reg _403470_403470 ; 
   reg __403470_403470;
   reg _403471_403471 ; 
   reg __403471_403471;
   reg _403472_403472 ; 
   reg __403472_403472;
   reg _403473_403473 ; 
   reg __403473_403473;
   reg _403474_403474 ; 
   reg __403474_403474;
   reg _403475_403475 ; 
   reg __403475_403475;
   reg _403476_403476 ; 
   reg __403476_403476;
   reg _403477_403477 ; 
   reg __403477_403477;
   reg _403478_403478 ; 
   reg __403478_403478;
   reg _403479_403479 ; 
   reg __403479_403479;
   reg _403480_403480 ; 
   reg __403480_403480;
   reg _403481_403481 ; 
   reg __403481_403481;
   reg _403482_403482 ; 
   reg __403482_403482;
   reg _403483_403483 ; 
   reg __403483_403483;
   reg _403484_403484 ; 
   reg __403484_403484;
   reg _403485_403485 ; 
   reg __403485_403485;
   reg _403486_403486 ; 
   reg __403486_403486;
   reg _403487_403487 ; 
   reg __403487_403487;
   reg _403488_403488 ; 
   reg __403488_403488;
   reg _403489_403489 ; 
   reg __403489_403489;
   reg _403490_403490 ; 
   reg __403490_403490;
   reg _403491_403491 ; 
   reg __403491_403491;
   reg _403492_403492 ; 
   reg __403492_403492;
   reg _403493_403493 ; 
   reg __403493_403493;
   reg _403494_403494 ; 
   reg __403494_403494;
   reg _403495_403495 ; 
   reg __403495_403495;
   reg _403496_403496 ; 
   reg __403496_403496;
   reg _403497_403497 ; 
   reg __403497_403497;
   reg _403498_403498 ; 
   reg __403498_403498;
   reg _403499_403499 ; 
   reg __403499_403499;
   reg _403500_403500 ; 
   reg __403500_403500;
   reg _403501_403501 ; 
   reg __403501_403501;
   reg _403502_403502 ; 
   reg __403502_403502;
   reg _403503_403503 ; 
   reg __403503_403503;
   reg _403504_403504 ; 
   reg __403504_403504;
   reg _403505_403505 ; 
   reg __403505_403505;
   reg _403506_403506 ; 
   reg __403506_403506;
   reg _403507_403507 ; 
   reg __403507_403507;
   reg _403508_403508 ; 
   reg __403508_403508;
   reg _403509_403509 ; 
   reg __403509_403509;
   reg _403510_403510 ; 
   reg __403510_403510;
   reg _403511_403511 ; 
   reg __403511_403511;
   reg _403512_403512 ; 
   reg __403512_403512;
   reg _403513_403513 ; 
   reg __403513_403513;
   reg _403514_403514 ; 
   reg __403514_403514;
   reg _403515_403515 ; 
   reg __403515_403515;
   reg _403516_403516 ; 
   reg __403516_403516;
   reg _403517_403517 ; 
   reg __403517_403517;
   reg _403518_403518 ; 
   reg __403518_403518;
   reg _403519_403519 ; 
   reg __403519_403519;
   reg _403520_403520 ; 
   reg __403520_403520;
   reg _403521_403521 ; 
   reg __403521_403521;
   reg _403522_403522 ; 
   reg __403522_403522;
   reg _403523_403523 ; 
   reg __403523_403523;
   reg _403524_403524 ; 
   reg __403524_403524;
   reg _403525_403525 ; 
   reg __403525_403525;
   reg _403526_403526 ; 
   reg __403526_403526;
   reg _403527_403527 ; 
   reg __403527_403527;
   reg _403528_403528 ; 
   reg __403528_403528;
   reg _403529_403529 ; 
   reg __403529_403529;
   reg _403530_403530 ; 
   reg __403530_403530;
   reg _403531_403531 ; 
   reg __403531_403531;
   reg _403532_403532 ; 
   reg __403532_403532;
   reg _403533_403533 ; 
   reg __403533_403533;
   reg _403534_403534 ; 
   reg __403534_403534;
   reg _403535_403535 ; 
   reg __403535_403535;
   reg _403536_403536 ; 
   reg __403536_403536;
   reg _403537_403537 ; 
   reg __403537_403537;
   reg _403538_403538 ; 
   reg __403538_403538;
   reg _403539_403539 ; 
   reg __403539_403539;
   reg _403540_403540 ; 
   reg __403540_403540;
   reg _403541_403541 ; 
   reg __403541_403541;
   reg _403542_403542 ; 
   reg __403542_403542;
   reg _403543_403543 ; 
   reg __403543_403543;
   reg _403544_403544 ; 
   reg __403544_403544;
   reg _403545_403545 ; 
   reg __403545_403545;
   reg _403546_403546 ; 
   reg __403546_403546;
   reg _403547_403547 ; 
   reg __403547_403547;
   reg _403548_403548 ; 
   reg __403548_403548;
   reg _403549_403549 ; 
   reg __403549_403549;
   reg _403550_403550 ; 
   reg __403550_403550;
   reg _403551_403551 ; 
   reg __403551_403551;
   reg _403552_403552 ; 
   reg __403552_403552;
   reg _403553_403553 ; 
   reg __403553_403553;
   reg _403554_403554 ; 
   reg __403554_403554;
   reg _403555_403555 ; 
   reg __403555_403555;
   reg _403556_403556 ; 
   reg __403556_403556;
   reg _403557_403557 ; 
   reg __403557_403557;
   reg _403558_403558 ; 
   reg __403558_403558;
   reg _403559_403559 ; 
   reg __403559_403559;
   reg _403560_403560 ; 
   reg __403560_403560;
   reg _403561_403561 ; 
   reg __403561_403561;
   reg _403562_403562 ; 
   reg __403562_403562;
   reg _403563_403563 ; 
   reg __403563_403563;
   reg _403564_403564 ; 
   reg __403564_403564;
   reg _403565_403565 ; 
   reg __403565_403565;
   reg _403566_403566 ; 
   reg __403566_403566;
   reg _403567_403567 ; 
   reg __403567_403567;
   reg _403568_403568 ; 
   reg __403568_403568;
   reg _403569_403569 ; 
   reg __403569_403569;
   reg _403570_403570 ; 
   reg __403570_403570;
   reg _403571_403571 ; 
   reg __403571_403571;
   reg _403572_403572 ; 
   reg __403572_403572;
   reg _403573_403573 ; 
   reg __403573_403573;
   reg _403574_403574 ; 
   reg __403574_403574;
   reg _403575_403575 ; 
   reg __403575_403575;
   reg _403576_403576 ; 
   reg __403576_403576;
   reg _403577_403577 ; 
   reg __403577_403577;
   reg _403578_403578 ; 
   reg __403578_403578;
   reg _403579_403579 ; 
   reg __403579_403579;
   reg _403580_403580 ; 
   reg __403580_403580;
   reg _403581_403581 ; 
   reg __403581_403581;
   reg _403582_403582 ; 
   reg __403582_403582;
   reg _403583_403583 ; 
   reg __403583_403583;
   reg _403584_403584 ; 
   reg __403584_403584;
   reg _403585_403585 ; 
   reg __403585_403585;
   reg _403586_403586 ; 
   reg __403586_403586;
   reg _403587_403587 ; 
   reg __403587_403587;
   reg _403588_403588 ; 
   reg __403588_403588;
   reg _403589_403589 ; 
   reg __403589_403589;
   reg _403590_403590 ; 
   reg __403590_403590;
   reg _403591_403591 ; 
   reg __403591_403591;
   reg _403592_403592 ; 
   reg __403592_403592;
   reg _403593_403593 ; 
   reg __403593_403593;
   reg _403594_403594 ; 
   reg __403594_403594;
   reg _403595_403595 ; 
   reg __403595_403595;
   reg _403596_403596 ; 
   reg __403596_403596;
   reg _403597_403597 ; 
   reg __403597_403597;
   reg _403598_403598 ; 
   reg __403598_403598;
   reg _403599_403599 ; 
   reg __403599_403599;
   reg _403600_403600 ; 
   reg __403600_403600;
   reg _403601_403601 ; 
   reg __403601_403601;
   reg _403602_403602 ; 
   reg __403602_403602;
   reg _403603_403603 ; 
   reg __403603_403603;
   reg _403604_403604 ; 
   reg __403604_403604;
   reg _403605_403605 ; 
   reg __403605_403605;
   reg _403606_403606 ; 
   reg __403606_403606;
   reg _403607_403607 ; 
   reg __403607_403607;
   reg _403608_403608 ; 
   reg __403608_403608;
   reg _403609_403609 ; 
   reg __403609_403609;
   reg _403610_403610 ; 
   reg __403610_403610;
   reg _403611_403611 ; 
   reg __403611_403611;
   reg _403612_403612 ; 
   reg __403612_403612;
   reg _403613_403613 ; 
   reg __403613_403613;
   reg _403614_403614 ; 
   reg __403614_403614;
   reg _403615_403615 ; 
   reg __403615_403615;
   reg _403616_403616 ; 
   reg __403616_403616;
   reg _403617_403617 ; 
   reg __403617_403617;
   reg _403618_403618 ; 
   reg __403618_403618;
   reg _403619_403619 ; 
   reg __403619_403619;
   reg _403620_403620 ; 
   reg __403620_403620;
   reg _403621_403621 ; 
   reg __403621_403621;
   reg _403622_403622 ; 
   reg __403622_403622;
   reg _403623_403623 ; 
   reg __403623_403623;
   reg _403624_403624 ; 
   reg __403624_403624;
   reg _403625_403625 ; 
   reg __403625_403625;
   reg _403626_403626 ; 
   reg __403626_403626;
   reg _403627_403627 ; 
   reg __403627_403627;
   reg _403628_403628 ; 
   reg __403628_403628;
   reg _403629_403629 ; 
   reg __403629_403629;
   reg _403630_403630 ; 
   reg __403630_403630;
   reg _403631_403631 ; 
   reg __403631_403631;
   reg _403632_403632 ; 
   reg __403632_403632;
   reg _403633_403633 ; 
   reg __403633_403633;
   reg _403634_403634 ; 
   reg __403634_403634;
   reg _403635_403635 ; 
   reg __403635_403635;
   reg _403636_403636 ; 
   reg __403636_403636;
   reg _403637_403637 ; 
   reg __403637_403637;
   reg _403638_403638 ; 
   reg __403638_403638;
   reg _403639_403639 ; 
   reg __403639_403639;
   reg _403640_403640 ; 
   reg __403640_403640;
   reg _403641_403641 ; 
   reg __403641_403641;
   reg _403642_403642 ; 
   reg __403642_403642;
   reg _403643_403643 ; 
   reg __403643_403643;
   reg _403644_403644 ; 
   reg __403644_403644;
   reg _403645_403645 ; 
   reg __403645_403645;
   reg _403646_403646 ; 
   reg __403646_403646;
   reg _403647_403647 ; 
   reg __403647_403647;
   reg _403648_403648 ; 
   reg __403648_403648;
   reg _403649_403649 ; 
   reg __403649_403649;
   reg _403650_403650 ; 
   reg __403650_403650;
   reg _403651_403651 ; 
   reg __403651_403651;
   reg _403652_403652 ; 
   reg __403652_403652;
   reg _403653_403653 ; 
   reg __403653_403653;
   reg _403654_403654 ; 
   reg __403654_403654;
   reg _403655_403655 ; 
   reg __403655_403655;
   reg _403656_403656 ; 
   reg __403656_403656;
   reg _403657_403657 ; 
   reg __403657_403657;
   reg _403658_403658 ; 
   reg __403658_403658;
   reg _403659_403659 ; 
   reg __403659_403659;
   reg _403660_403660 ; 
   reg __403660_403660;
   reg _403661_403661 ; 
   reg __403661_403661;
   reg _403662_403662 ; 
   reg __403662_403662;
   reg _403663_403663 ; 
   reg __403663_403663;
   reg _403664_403664 ; 
   reg __403664_403664;
   reg _403665_403665 ; 
   reg __403665_403665;
   reg _403666_403666 ; 
   reg __403666_403666;
   reg _403667_403667 ; 
   reg __403667_403667;
   reg _403668_403668 ; 
   reg __403668_403668;
   reg _403669_403669 ; 
   reg __403669_403669;
   reg _403670_403670 ; 
   reg __403670_403670;
   reg _403671_403671 ; 
   reg __403671_403671;
   reg _403672_403672 ; 
   reg __403672_403672;
   reg _403673_403673 ; 
   reg __403673_403673;
   reg _403674_403674 ; 
   reg __403674_403674;
   reg _403675_403675 ; 
   reg __403675_403675;
   reg _403676_403676 ; 
   reg __403676_403676;
   reg _403677_403677 ; 
   reg __403677_403677;
   reg _403678_403678 ; 
   reg __403678_403678;
   reg _403679_403679 ; 
   reg __403679_403679;
   reg _403680_403680 ; 
   reg __403680_403680;
   reg _403681_403681 ; 
   reg __403681_403681;
   reg _403682_403682 ; 
   reg __403682_403682;
   reg _403683_403683 ; 
   reg __403683_403683;
   reg _403684_403684 ; 
   reg __403684_403684;
   reg _403685_403685 ; 
   reg __403685_403685;
   reg _403686_403686 ; 
   reg __403686_403686;
   reg _403687_403687 ; 
   reg __403687_403687;
   reg _403688_403688 ; 
   reg __403688_403688;
   reg _403689_403689 ; 
   reg __403689_403689;
   reg _403690_403690 ; 
   reg __403690_403690;
   reg _403691_403691 ; 
   reg __403691_403691;
   reg _403692_403692 ; 
   reg __403692_403692;
   reg _403693_403693 ; 
   reg __403693_403693;
   reg _403694_403694 ; 
   reg __403694_403694;
   reg _403695_403695 ; 
   reg __403695_403695;
   reg _403696_403696 ; 
   reg __403696_403696;
   reg _403697_403697 ; 
   reg __403697_403697;
   reg _403698_403698 ; 
   reg __403698_403698;
   reg _403699_403699 ; 
   reg __403699_403699;
   reg _403700_403700 ; 
   reg __403700_403700;
   reg _403701_403701 ; 
   reg __403701_403701;
   reg _403702_403702 ; 
   reg __403702_403702;
   reg _403703_403703 ; 
   reg __403703_403703;
   reg _403704_403704 ; 
   reg __403704_403704;
   reg _403705_403705 ; 
   reg __403705_403705;
   reg _403706_403706 ; 
   reg __403706_403706;
   reg _403707_403707 ; 
   reg __403707_403707;
   reg _403708_403708 ; 
   reg __403708_403708;
   reg _403709_403709 ; 
   reg __403709_403709;
   reg _403710_403710 ; 
   reg __403710_403710;
   reg _403711_403711 ; 
   reg __403711_403711;
   reg _403712_403712 ; 
   reg __403712_403712;
   reg _403713_403713 ; 
   reg __403713_403713;
   reg _403714_403714 ; 
   reg __403714_403714;
   reg _403715_403715 ; 
   reg __403715_403715;
   reg _403716_403716 ; 
   reg __403716_403716;
   reg _403717_403717 ; 
   reg __403717_403717;
   reg _403718_403718 ; 
   reg __403718_403718;
   reg _403719_403719 ; 
   reg __403719_403719;
   reg _403720_403720 ; 
   reg __403720_403720;
   reg _403721_403721 ; 
   reg __403721_403721;
   reg _403722_403722 ; 
   reg __403722_403722;
   reg _403723_403723 ; 
   reg __403723_403723;
   reg _403724_403724 ; 
   reg __403724_403724;
   reg _403725_403725 ; 
   reg __403725_403725;
   reg _403726_403726 ; 
   reg __403726_403726;
   reg _403727_403727 ; 
   reg __403727_403727;
   reg _403728_403728 ; 
   reg __403728_403728;
   reg _403729_403729 ; 
   reg __403729_403729;
   reg _403730_403730 ; 
   reg __403730_403730;
   reg _403731_403731 ; 
   reg __403731_403731;
   reg _403732_403732 ; 
   reg __403732_403732;
   reg _403733_403733 ; 
   reg __403733_403733;
   reg _403734_403734 ; 
   reg __403734_403734;
   reg _403735_403735 ; 
   reg __403735_403735;
   reg _403736_403736 ; 
   reg __403736_403736;
   reg _403737_403737 ; 
   reg __403737_403737;
   reg _403738_403738 ; 
   reg __403738_403738;
   reg _403739_403739 ; 
   reg __403739_403739;
   reg _403740_403740 ; 
   reg __403740_403740;
   reg _403741_403741 ; 
   reg __403741_403741;
   reg _403742_403742 ; 
   reg __403742_403742;
   reg _403743_403743 ; 
   reg __403743_403743;
   reg _403744_403744 ; 
   reg __403744_403744;
   reg _403745_403745 ; 
   reg __403745_403745;
   reg _403746_403746 ; 
   reg __403746_403746;
   reg _403747_403747 ; 
   reg __403747_403747;
   reg _403748_403748 ; 
   reg __403748_403748;
   reg _403749_403749 ; 
   reg __403749_403749;
   reg _403750_403750 ; 
   reg __403750_403750;
   reg _403751_403751 ; 
   reg __403751_403751;
   reg _403752_403752 ; 
   reg __403752_403752;
   reg _403753_403753 ; 
   reg __403753_403753;
   reg _403754_403754 ; 
   reg __403754_403754;
   reg _403755_403755 ; 
   reg __403755_403755;
   reg _403756_403756 ; 
   reg __403756_403756;
   reg _403757_403757 ; 
   reg __403757_403757;
   reg _403758_403758 ; 
   reg __403758_403758;
   reg _403759_403759 ; 
   reg __403759_403759;
   reg _403760_403760 ; 
   reg __403760_403760;
   reg _403761_403761 ; 
   reg __403761_403761;
   reg _403762_403762 ; 
   reg __403762_403762;
   reg _403763_403763 ; 
   reg __403763_403763;
   reg _403764_403764 ; 
   reg __403764_403764;
   reg _403765_403765 ; 
   reg __403765_403765;
   reg _403766_403766 ; 
   reg __403766_403766;
   reg _403767_403767 ; 
   reg __403767_403767;
   reg _403768_403768 ; 
   reg __403768_403768;
   reg _403769_403769 ; 
   reg __403769_403769;
   reg _403770_403770 ; 
   reg __403770_403770;
   reg _403771_403771 ; 
   reg __403771_403771;
   reg _403772_403772 ; 
   reg __403772_403772;
   reg _403773_403773 ; 
   reg __403773_403773;
   reg _403774_403774 ; 
   reg __403774_403774;
   reg _403775_403775 ; 
   reg __403775_403775;
   reg _403776_403776 ; 
   reg __403776_403776;
   reg _403777_403777 ; 
   reg __403777_403777;
   reg _403778_403778 ; 
   reg __403778_403778;
   reg _403779_403779 ; 
   reg __403779_403779;
   reg _403780_403780 ; 
   reg __403780_403780;
   reg _403781_403781 ; 
   reg __403781_403781;
   reg _403782_403782 ; 
   reg __403782_403782;
   reg _403783_403783 ; 
   reg __403783_403783;
   reg _403784_403784 ; 
   reg __403784_403784;
   reg _403785_403785 ; 
   reg __403785_403785;
   reg _403786_403786 ; 
   reg __403786_403786;
   reg _403787_403787 ; 
   reg __403787_403787;
   reg _403788_403788 ; 
   reg __403788_403788;
   reg _403789_403789 ; 
   reg __403789_403789;
   reg _403790_403790 ; 
   reg __403790_403790;
   reg _403791_403791 ; 
   reg __403791_403791;
   reg _403792_403792 ; 
   reg __403792_403792;
   reg _403793_403793 ; 
   reg __403793_403793;
   reg _403794_403794 ; 
   reg __403794_403794;
   reg _403795_403795 ; 
   reg __403795_403795;
   reg _403796_403796 ; 
   reg __403796_403796;
   reg _403797_403797 ; 
   reg __403797_403797;
   reg _403798_403798 ; 
   reg __403798_403798;
   reg _403799_403799 ; 
   reg __403799_403799;
   reg _403800_403800 ; 
   reg __403800_403800;
   reg _403801_403801 ; 
   reg __403801_403801;
   reg _403802_403802 ; 
   reg __403802_403802;
   reg _403803_403803 ; 
   reg __403803_403803;
   reg _403804_403804 ; 
   reg __403804_403804;
   reg _403805_403805 ; 
   reg __403805_403805;
   reg _403806_403806 ; 
   reg __403806_403806;
   reg _403807_403807 ; 
   reg __403807_403807;
   reg _403808_403808 ; 
   reg __403808_403808;
   reg _403809_403809 ; 
   reg __403809_403809;
   reg _403810_403810 ; 
   reg __403810_403810;
   reg _403811_403811 ; 
   reg __403811_403811;
   reg _403812_403812 ; 
   reg __403812_403812;
   reg _403813_403813 ; 
   reg __403813_403813;
   reg _403814_403814 ; 
   reg __403814_403814;
   reg _403815_403815 ; 
   reg __403815_403815;
   reg _403816_403816 ; 
   reg __403816_403816;
   reg _403817_403817 ; 
   reg __403817_403817;
   reg _403818_403818 ; 
   reg __403818_403818;
   reg _403819_403819 ; 
   reg __403819_403819;
   reg _403820_403820 ; 
   reg __403820_403820;
   reg _403821_403821 ; 
   reg __403821_403821;
   reg _403822_403822 ; 
   reg __403822_403822;
   reg _403823_403823 ; 
   reg __403823_403823;
   reg _403824_403824 ; 
   reg __403824_403824;
   reg _403825_403825 ; 
   reg __403825_403825;
   reg _403826_403826 ; 
   reg __403826_403826;
   reg _403827_403827 ; 
   reg __403827_403827;
   reg _403828_403828 ; 
   reg __403828_403828;
   reg _403829_403829 ; 
   reg __403829_403829;
   reg _403830_403830 ; 
   reg __403830_403830;
   reg _403831_403831 ; 
   reg __403831_403831;
   reg _403832_403832 ; 
   reg __403832_403832;
   reg _403833_403833 ; 
   reg __403833_403833;
   reg _403834_403834 ; 
   reg __403834_403834;
   reg _403835_403835 ; 
   reg __403835_403835;
   reg _403836_403836 ; 
   reg __403836_403836;
   reg _403837_403837 ; 
   reg __403837_403837;
   reg _403838_403838 ; 
   reg __403838_403838;
   reg _403839_403839 ; 
   reg __403839_403839;
   reg _403840_403840 ; 
   reg __403840_403840;
   reg _403841_403841 ; 
   reg __403841_403841;
   reg _403842_403842 ; 
   reg __403842_403842;
   reg _403843_403843 ; 
   reg __403843_403843;
   reg _403844_403844 ; 
   reg __403844_403844;
   reg _403845_403845 ; 
   reg __403845_403845;
   reg _403846_403846 ; 
   reg __403846_403846;
   reg _403847_403847 ; 
   reg __403847_403847;
   reg _403848_403848 ; 
   reg __403848_403848;
   reg _403849_403849 ; 
   reg __403849_403849;
   reg _403850_403850 ; 
   reg __403850_403850;
   reg _403851_403851 ; 
   reg __403851_403851;
   reg _403852_403852 ; 
   reg __403852_403852;
   reg _403853_403853 ; 
   reg __403853_403853;
   reg _403854_403854 ; 
   reg __403854_403854;
   reg _403855_403855 ; 
   reg __403855_403855;
   reg _403856_403856 ; 
   reg __403856_403856;
   reg _403857_403857 ; 
   reg __403857_403857;
   reg _403858_403858 ; 
   reg __403858_403858;
   reg _403859_403859 ; 
   reg __403859_403859;
   reg _403860_403860 ; 
   reg __403860_403860;
   reg _403861_403861 ; 
   reg __403861_403861;
   reg _403862_403862 ; 
   reg __403862_403862;
   reg _403863_403863 ; 
   reg __403863_403863;
   reg _403864_403864 ; 
   reg __403864_403864;
   reg _403865_403865 ; 
   reg __403865_403865;
   reg _403866_403866 ; 
   reg __403866_403866;
   reg _403867_403867 ; 
   reg __403867_403867;
   reg _403868_403868 ; 
   reg __403868_403868;
   reg _403869_403869 ; 
   reg __403869_403869;
   reg _403870_403870 ; 
   reg __403870_403870;
   reg _403871_403871 ; 
   reg __403871_403871;
   reg _403872_403872 ; 
   reg __403872_403872;
   reg _403873_403873 ; 
   reg __403873_403873;
   reg _403874_403874 ; 
   reg __403874_403874;
   reg _403875_403875 ; 
   reg __403875_403875;
   reg _403876_403876 ; 
   reg __403876_403876;
   reg _403877_403877 ; 
   reg __403877_403877;
   reg _403878_403878 ; 
   reg __403878_403878;
   reg _403879_403879 ; 
   reg __403879_403879;
   reg _403880_403880 ; 
   reg __403880_403880;
   reg _403881_403881 ; 
   reg __403881_403881;
   reg _403882_403882 ; 
   reg __403882_403882;
   reg _403883_403883 ; 
   reg __403883_403883;
   reg _403884_403884 ; 
   reg __403884_403884;
   reg _403885_403885 ; 
   reg __403885_403885;
   reg _403886_403886 ; 
   reg __403886_403886;
   reg _403887_403887 ; 
   reg __403887_403887;
   reg _403888_403888 ; 
   reg __403888_403888;
   reg _403889_403889 ; 
   reg __403889_403889;
   reg _403890_403890 ; 
   reg __403890_403890;
   reg _403891_403891 ; 
   reg __403891_403891;
   reg _403892_403892 ; 
   reg __403892_403892;
   reg _403893_403893 ; 
   reg __403893_403893;
   reg _403894_403894 ; 
   reg __403894_403894;
   reg _403895_403895 ; 
   reg __403895_403895;
   reg _403896_403896 ; 
   reg __403896_403896;
   reg _403897_403897 ; 
   reg __403897_403897;
   reg _403898_403898 ; 
   reg __403898_403898;
   reg _403899_403899 ; 
   reg __403899_403899;
   reg _403900_403900 ; 
   reg __403900_403900;
   reg _403901_403901 ; 
   reg __403901_403901;
   reg _403902_403902 ; 
   reg __403902_403902;
   reg _403903_403903 ; 
   reg __403903_403903;
   reg _403904_403904 ; 
   reg __403904_403904;
   reg _403905_403905 ; 
   reg __403905_403905;
   reg _403906_403906 ; 
   reg __403906_403906;
   reg _403907_403907 ; 
   reg __403907_403907;
   reg _403908_403908 ; 
   reg __403908_403908;
   reg _403909_403909 ; 
   reg __403909_403909;
   reg _403910_403910 ; 
   reg __403910_403910;
   reg _403911_403911 ; 
   reg __403911_403911;
   reg _403912_403912 ; 
   reg __403912_403912;
   reg _403913_403913 ; 
   reg __403913_403913;
   reg _403914_403914 ; 
   reg __403914_403914;
   reg _403915_403915 ; 
   reg __403915_403915;
   reg _403916_403916 ; 
   reg __403916_403916;
   reg _403917_403917 ; 
   reg __403917_403917;
   reg _403918_403918 ; 
   reg __403918_403918;
   reg _403919_403919 ; 
   reg __403919_403919;
   reg _403920_403920 ; 
   reg __403920_403920;
   reg _403921_403921 ; 
   reg __403921_403921;
   reg _403922_403922 ; 
   reg __403922_403922;
   reg _403923_403923 ; 
   reg __403923_403923;
   reg _403924_403924 ; 
   reg __403924_403924;
   reg _403925_403925 ; 
   reg __403925_403925;
   reg _403926_403926 ; 
   reg __403926_403926;
   reg _403927_403927 ; 
   reg __403927_403927;
   reg _403928_403928 ; 
   reg __403928_403928;
   reg _403929_403929 ; 
   reg __403929_403929;
   reg _403930_403930 ; 
   reg __403930_403930;
   reg _403931_403931 ; 
   reg __403931_403931;
   reg _403932_403932 ; 
   reg __403932_403932;
   reg _403933_403933 ; 
   reg __403933_403933;
   reg _403934_403934 ; 
   reg __403934_403934;
   reg _403935_403935 ; 
   reg __403935_403935;
   reg _403936_403936 ; 
   reg __403936_403936;
   reg _403937_403937 ; 
   reg __403937_403937;
   reg _403938_403938 ; 
   reg __403938_403938;
   reg _403939_403939 ; 
   reg __403939_403939;
   reg _403940_403940 ; 
   reg __403940_403940;
   reg _403941_403941 ; 
   reg __403941_403941;
   reg _403942_403942 ; 
   reg __403942_403942;
   reg _403943_403943 ; 
   reg __403943_403943;
   reg _403944_403944 ; 
   reg __403944_403944;
   reg _403945_403945 ; 
   reg __403945_403945;
   reg _403946_403946 ; 
   reg __403946_403946;
   reg _403947_403947 ; 
   reg __403947_403947;
   reg _403948_403948 ; 
   reg __403948_403948;
   reg _403949_403949 ; 
   reg __403949_403949;
   reg _403950_403950 ; 
   reg __403950_403950;
   reg _403951_403951 ; 
   reg __403951_403951;
   reg _403952_403952 ; 
   reg __403952_403952;
   reg _403953_403953 ; 
   reg __403953_403953;
   reg _403954_403954 ; 
   reg __403954_403954;
   reg _403955_403955 ; 
   reg __403955_403955;
   reg _403956_403956 ; 
   reg __403956_403956;
   reg _403957_403957 ; 
   reg __403957_403957;
   reg _403958_403958 ; 
   reg __403958_403958;
   reg _403959_403959 ; 
   reg __403959_403959;
   reg _403960_403960 ; 
   reg __403960_403960;
   reg _403961_403961 ; 
   reg __403961_403961;
   reg _403962_403962 ; 
   reg __403962_403962;
   reg _403963_403963 ; 
   reg __403963_403963;
   reg _403964_403964 ; 
   reg __403964_403964;
   reg _403965_403965 ; 
   reg __403965_403965;
   reg _403966_403966 ; 
   reg __403966_403966;
   reg _403967_403967 ; 
   reg __403967_403967;
   reg _403968_403968 ; 
   reg __403968_403968;
   reg _403969_403969 ; 
   reg __403969_403969;
   reg _403970_403970 ; 
   reg __403970_403970;
   reg _403971_403971 ; 
   reg __403971_403971;
   reg _403972_403972 ; 
   reg __403972_403972;
   reg _403973_403973 ; 
   reg __403973_403973;
   reg _403974_403974 ; 
   reg __403974_403974;
   reg _403975_403975 ; 
   reg __403975_403975;
   reg _403976_403976 ; 
   reg __403976_403976;
   reg _403977_403977 ; 
   reg __403977_403977;
   reg _403978_403978 ; 
   reg __403978_403978;
   reg _403979_403979 ; 
   reg __403979_403979;
   reg _403980_403980 ; 
   reg __403980_403980;
   reg _403981_403981 ; 
   reg __403981_403981;
   reg _403982_403982 ; 
   reg __403982_403982;
   reg _403983_403983 ; 
   reg __403983_403983;
   reg _403984_403984 ; 
   reg __403984_403984;
   reg _403985_403985 ; 
   reg __403985_403985;
   reg _403986_403986 ; 
   reg __403986_403986;
   reg _403987_403987 ; 
   reg __403987_403987;
   reg _403988_403988 ; 
   reg __403988_403988;
   reg _403989_403989 ; 
   reg __403989_403989;
   reg _403990_403990 ; 
   reg __403990_403990;
   reg _403991_403991 ; 
   reg __403991_403991;
   reg _403992_403992 ; 
   reg __403992_403992;
   reg _403993_403993 ; 
   reg __403993_403993;
   reg _403994_403994 ; 
   reg __403994_403994;
   reg _403995_403995 ; 
   reg __403995_403995;
   reg _403996_403996 ; 
   reg __403996_403996;
   reg _403997_403997 ; 
   reg __403997_403997;
   reg _403998_403998 ; 
   reg __403998_403998;
   reg _403999_403999 ; 
   reg __403999_403999;
   reg _404000_404000 ; 
   reg __404000_404000;
   reg _404001_404001 ; 
   reg __404001_404001;
   reg _404002_404002 ; 
   reg __404002_404002;
   reg _404003_404003 ; 
   reg __404003_404003;
   reg _404004_404004 ; 
   reg __404004_404004;
   reg _404005_404005 ; 
   reg __404005_404005;
   reg _404006_404006 ; 
   reg __404006_404006;
   reg _404007_404007 ; 
   reg __404007_404007;
   reg _404008_404008 ; 
   reg __404008_404008;
   reg _404009_404009 ; 
   reg __404009_404009;
   reg _404010_404010 ; 
   reg __404010_404010;
   reg _404011_404011 ; 
   reg __404011_404011;
   reg _404012_404012 ; 
   reg __404012_404012;
   reg _404013_404013 ; 
   reg __404013_404013;
   reg _404014_404014 ; 
   reg __404014_404014;
   reg _404015_404015 ; 
   reg __404015_404015;
   reg _404016_404016 ; 
   reg __404016_404016;
   reg _404017_404017 ; 
   reg __404017_404017;
   reg _404018_404018 ; 
   reg __404018_404018;
   reg _404019_404019 ; 
   reg __404019_404019;
   reg _404020_404020 ; 
   reg __404020_404020;
   reg _404021_404021 ; 
   reg __404021_404021;
   reg _404022_404022 ; 
   reg __404022_404022;
   reg _404023_404023 ; 
   reg __404023_404023;
   reg _404024_404024 ; 
   reg __404024_404024;
   reg _404025_404025 ; 
   reg __404025_404025;
   reg _404026_404026 ; 
   reg __404026_404026;
   reg _404027_404027 ; 
   reg __404027_404027;
   reg _404028_404028 ; 
   reg __404028_404028;
   reg _404029_404029 ; 
   reg __404029_404029;
   reg _404030_404030 ; 
   reg __404030_404030;
   reg _404031_404031 ; 
   reg __404031_404031;
   reg _404032_404032 ; 
   reg __404032_404032;
   reg _404033_404033 ; 
   reg __404033_404033;
   reg _404034_404034 ; 
   reg __404034_404034;
   reg _404035_404035 ; 
   reg __404035_404035;
   reg _404036_404036 ; 
   reg __404036_404036;
   reg _404037_404037 ; 
   reg __404037_404037;
   reg _404038_404038 ; 
   reg __404038_404038;
   reg _404039_404039 ; 
   reg __404039_404039;
   reg _404040_404040 ; 
   reg __404040_404040;
   reg _404041_404041 ; 
   reg __404041_404041;
   reg _404042_404042 ; 
   reg __404042_404042;
   reg _404043_404043 ; 
   reg __404043_404043;
   reg _404044_404044 ; 
   reg __404044_404044;
   reg _404045_404045 ; 
   reg __404045_404045;
   reg _404046_404046 ; 
   reg __404046_404046;
   reg _404047_404047 ; 
   reg __404047_404047;
   reg _404048_404048 ; 
   reg __404048_404048;
   reg _404049_404049 ; 
   reg __404049_404049;
   reg _404050_404050 ; 
   reg __404050_404050;
   reg _404051_404051 ; 
   reg __404051_404051;
   reg _404052_404052 ; 
   reg __404052_404052;
   reg _404053_404053 ; 
   reg __404053_404053;
   reg _404054_404054 ; 
   reg __404054_404054;
   reg _404055_404055 ; 
   reg __404055_404055;
   reg _404056_404056 ; 
   reg __404056_404056;
   reg _404057_404057 ; 
   reg __404057_404057;
   reg _404058_404058 ; 
   reg __404058_404058;
   reg _404059_404059 ; 
   reg __404059_404059;
   reg _404060_404060 ; 
   reg __404060_404060;
   reg _404061_404061 ; 
   reg __404061_404061;
   reg _404062_404062 ; 
   reg __404062_404062;
   reg _404063_404063 ; 
   reg __404063_404063;
   reg _404064_404064 ; 
   reg __404064_404064;
   reg _404065_404065 ; 
   reg __404065_404065;
   reg _404066_404066 ; 
   reg __404066_404066;
   reg _404067_404067 ; 
   reg __404067_404067;
   reg _404068_404068 ; 
   reg __404068_404068;
   reg _404069_404069 ; 
   reg __404069_404069;
   reg _404070_404070 ; 
   reg __404070_404070;
   reg _404071_404071 ; 
   reg __404071_404071;
   reg _404072_404072 ; 
   reg __404072_404072;
   reg _404073_404073 ; 
   reg __404073_404073;
   reg _404074_404074 ; 
   reg __404074_404074;
   reg _404075_404075 ; 
   reg __404075_404075;
   reg _404076_404076 ; 
   reg __404076_404076;
   reg _404077_404077 ; 
   reg __404077_404077;
   reg _404078_404078 ; 
   reg __404078_404078;
   reg _404079_404079 ; 
   reg __404079_404079;
   reg _404080_404080 ; 
   reg __404080_404080;
   reg _404081_404081 ; 
   reg __404081_404081;
   reg _404082_404082 ; 
   reg __404082_404082;
   reg _404083_404083 ; 
   reg __404083_404083;
   reg _404084_404084 ; 
   reg __404084_404084;
   reg _404085_404085 ; 
   reg __404085_404085;
   reg _404086_404086 ; 
   reg __404086_404086;
   reg _404087_404087 ; 
   reg __404087_404087;
   reg _404088_404088 ; 
   reg __404088_404088;
   reg _404089_404089 ; 
   reg __404089_404089;
   reg _404090_404090 ; 
   reg __404090_404090;
   reg _404091_404091 ; 
   reg __404091_404091;
   reg _404092_404092 ; 
   reg __404092_404092;
   reg _404093_404093 ; 
   reg __404093_404093;
   reg _404094_404094 ; 
   reg __404094_404094;
   reg _404095_404095 ; 
   reg __404095_404095;
   reg _404096_404096 ; 
   reg __404096_404096;
   reg _404097_404097 ; 
   reg __404097_404097;
   reg _404098_404098 ; 
   reg __404098_404098;
   reg _404099_404099 ; 
   reg __404099_404099;
   reg _404100_404100 ; 
   reg __404100_404100;
   reg _404101_404101 ; 
   reg __404101_404101;
   reg _404102_404102 ; 
   reg __404102_404102;
   reg _404103_404103 ; 
   reg __404103_404103;
   reg _404104_404104 ; 
   reg __404104_404104;
   reg _404105_404105 ; 
   reg __404105_404105;
   reg _404106_404106 ; 
   reg __404106_404106;
   reg _404107_404107 ; 
   reg __404107_404107;
   reg _404108_404108 ; 
   reg __404108_404108;
   reg _404109_404109 ; 
   reg __404109_404109;
   reg _404110_404110 ; 
   reg __404110_404110;
   reg _404111_404111 ; 
   reg __404111_404111;
   reg _404112_404112 ; 
   reg __404112_404112;
   reg _404113_404113 ; 
   reg __404113_404113;
   reg _404114_404114 ; 
   reg __404114_404114;
   reg _404115_404115 ; 
   reg __404115_404115;
   reg _404116_404116 ; 
   reg __404116_404116;
   reg _404117_404117 ; 
   reg __404117_404117;
   reg _404118_404118 ; 
   reg __404118_404118;
   reg _404119_404119 ; 
   reg __404119_404119;
   reg _404120_404120 ; 
   reg __404120_404120;
   reg _404121_404121 ; 
   reg __404121_404121;
   reg _404122_404122 ; 
   reg __404122_404122;
   reg _404123_404123 ; 
   reg __404123_404123;
   reg _404124_404124 ; 
   reg __404124_404124;
   reg _404125_404125 ; 
   reg __404125_404125;
   reg _404126_404126 ; 
   reg __404126_404126;
   reg _404127_404127 ; 
   reg __404127_404127;
   reg _404128_404128 ; 
   reg __404128_404128;
   reg _404129_404129 ; 
   reg __404129_404129;
   reg _404130_404130 ; 
   reg __404130_404130;
   reg _404131_404131 ; 
   reg __404131_404131;
   reg _404132_404132 ; 
   reg __404132_404132;
   reg _404133_404133 ; 
   reg __404133_404133;
   reg _404134_404134 ; 
   reg __404134_404134;
   reg _404135_404135 ; 
   reg __404135_404135;
   reg _404136_404136 ; 
   reg __404136_404136;
   reg _404137_404137 ; 
   reg __404137_404137;
   reg _404138_404138 ; 
   reg __404138_404138;
   reg _404139_404139 ; 
   reg __404139_404139;
   reg _404140_404140 ; 
   reg __404140_404140;
   reg _404141_404141 ; 
   reg __404141_404141;
   reg _404142_404142 ; 
   reg __404142_404142;
   reg _404143_404143 ; 
   reg __404143_404143;
   reg _404144_404144 ; 
   reg __404144_404144;
   reg _404145_404145 ; 
   reg __404145_404145;
   reg _404146_404146 ; 
   reg __404146_404146;
   reg _404147_404147 ; 
   reg __404147_404147;
   reg _404148_404148 ; 
   reg __404148_404148;
   reg _404149_404149 ; 
   reg __404149_404149;
   reg _404150_404150 ; 
   reg __404150_404150;
   reg _404151_404151 ; 
   reg __404151_404151;
   reg _404152_404152 ; 
   reg __404152_404152;
   reg _404153_404153 ; 
   reg __404153_404153;
   reg _404154_404154 ; 
   reg __404154_404154;
   reg _404155_404155 ; 
   reg __404155_404155;
   reg _404156_404156 ; 
   reg __404156_404156;
   reg _404157_404157 ; 
   reg __404157_404157;
   reg _404158_404158 ; 
   reg __404158_404158;
   reg _404159_404159 ; 
   reg __404159_404159;
   reg _404160_404160 ; 
   reg __404160_404160;
   reg _404161_404161 ; 
   reg __404161_404161;
   reg _404162_404162 ; 
   reg __404162_404162;
   reg _404163_404163 ; 
   reg __404163_404163;
   reg _404164_404164 ; 
   reg __404164_404164;
   reg _404165_404165 ; 
   reg __404165_404165;
   reg _404166_404166 ; 
   reg __404166_404166;
   reg _404167_404167 ; 
   reg __404167_404167;
   reg _404168_404168 ; 
   reg __404168_404168;
   reg _404169_404169 ; 
   reg __404169_404169;
   reg _404170_404170 ; 
   reg __404170_404170;
   reg _404171_404171 ; 
   reg __404171_404171;
   reg _404172_404172 ; 
   reg __404172_404172;
   reg _404173_404173 ; 
   reg __404173_404173;
   reg _404174_404174 ; 
   reg __404174_404174;
   reg _404175_404175 ; 
   reg __404175_404175;
   reg _404176_404176 ; 
   reg __404176_404176;
   reg _404177_404177 ; 
   reg __404177_404177;
   reg _404178_404178 ; 
   reg __404178_404178;
   reg _404179_404179 ; 
   reg __404179_404179;
   reg _404180_404180 ; 
   reg __404180_404180;
   reg _404181_404181 ; 
   reg __404181_404181;
   reg _404182_404182 ; 
   reg __404182_404182;
   reg _404183_404183 ; 
   reg __404183_404183;
   reg _404184_404184 ; 
   reg __404184_404184;
   reg _404185_404185 ; 
   reg __404185_404185;
   reg _404186_404186 ; 
   reg __404186_404186;
   reg _404187_404187 ; 
   reg __404187_404187;
   reg _404188_404188 ; 
   reg __404188_404188;
   reg _404189_404189 ; 
   reg __404189_404189;
   reg _404190_404190 ; 
   reg __404190_404190;
   reg _404191_404191 ; 
   reg __404191_404191;
   reg _404192_404192 ; 
   reg __404192_404192;
   reg _404193_404193 ; 
   reg __404193_404193;
   reg _404194_404194 ; 
   reg __404194_404194;
   reg _404195_404195 ; 
   reg __404195_404195;
   reg _404196_404196 ; 
   reg __404196_404196;
   reg _404197_404197 ; 
   reg __404197_404197;
   reg _404198_404198 ; 
   reg __404198_404198;
   reg _404199_404199 ; 
   reg __404199_404199;
   reg _404200_404200 ; 
   reg __404200_404200;
   reg _404201_404201 ; 
   reg __404201_404201;
   reg _404202_404202 ; 
   reg __404202_404202;
   reg _404203_404203 ; 
   reg __404203_404203;
   reg _404204_404204 ; 
   reg __404204_404204;
   reg _404205_404205 ; 
   reg __404205_404205;
   reg _404206_404206 ; 
   reg __404206_404206;
   reg _404207_404207 ; 
   reg __404207_404207;
   reg _404208_404208 ; 
   reg __404208_404208;
   reg _404209_404209 ; 
   reg __404209_404209;
   reg _404210_404210 ; 
   reg __404210_404210;
   reg _404211_404211 ; 
   reg __404211_404211;
   reg _404212_404212 ; 
   reg __404212_404212;
   reg _404213_404213 ; 
   reg __404213_404213;
   reg _404214_404214 ; 
   reg __404214_404214;
   reg _404215_404215 ; 
   reg __404215_404215;
   reg _404216_404216 ; 
   reg __404216_404216;
   reg _404217_404217 ; 
   reg __404217_404217;
   reg _404218_404218 ; 
   reg __404218_404218;
   reg _404219_404219 ; 
   reg __404219_404219;
   reg _404220_404220 ; 
   reg __404220_404220;
   reg _404221_404221 ; 
   reg __404221_404221;
   reg _404222_404222 ; 
   reg __404222_404222;
   reg _404223_404223 ; 
   reg __404223_404223;
   reg _404224_404224 ; 
   reg __404224_404224;
   reg _404225_404225 ; 
   reg __404225_404225;
   reg _404226_404226 ; 
   reg __404226_404226;
   reg _404227_404227 ; 
   reg __404227_404227;
   reg _404228_404228 ; 
   reg __404228_404228;
   reg _404229_404229 ; 
   reg __404229_404229;
   reg _404230_404230 ; 
   reg __404230_404230;
   reg _404231_404231 ; 
   reg __404231_404231;
   reg _404232_404232 ; 
   reg __404232_404232;
   reg _404233_404233 ; 
   reg __404233_404233;
   reg _404234_404234 ; 
   reg __404234_404234;
   reg _404235_404235 ; 
   reg __404235_404235;
   reg _404236_404236 ; 
   reg __404236_404236;
   reg _404237_404237 ; 
   reg __404237_404237;
   reg _404238_404238 ; 
   reg __404238_404238;
   reg _404239_404239 ; 
   reg __404239_404239;
   reg _404240_404240 ; 
   reg __404240_404240;
   reg _404241_404241 ; 
   reg __404241_404241;
   reg _404242_404242 ; 
   reg __404242_404242;
   reg _404243_404243 ; 
   reg __404243_404243;
   reg _404244_404244 ; 
   reg __404244_404244;
   reg _404245_404245 ; 
   reg __404245_404245;
   reg _404246_404246 ; 
   reg __404246_404246;
   reg _404247_404247 ; 
   reg __404247_404247;
   reg _404248_404248 ; 
   reg __404248_404248;
   reg _404249_404249 ; 
   reg __404249_404249;
   reg _404250_404250 ; 
   reg __404250_404250;
   reg _404251_404251 ; 
   reg __404251_404251;
   reg _404252_404252 ; 
   reg __404252_404252;
   reg _404253_404253 ; 
   reg __404253_404253;
   reg _404254_404254 ; 
   reg __404254_404254;
   reg _404255_404255 ; 
   reg __404255_404255;
   reg _404256_404256 ; 
   reg __404256_404256;
   reg _404257_404257 ; 
   reg __404257_404257;
   reg _404258_404258 ; 
   reg __404258_404258;
   reg _404259_404259 ; 
   reg __404259_404259;
   reg _404260_404260 ; 
   reg __404260_404260;
   reg _404261_404261 ; 
   reg __404261_404261;
   reg _404262_404262 ; 
   reg __404262_404262;
   reg _404263_404263 ; 
   reg __404263_404263;
   reg _404264_404264 ; 
   reg __404264_404264;
   reg _404265_404265 ; 
   reg __404265_404265;
   reg _404266_404266 ; 
   reg __404266_404266;
   reg _404267_404267 ; 
   reg __404267_404267;
   reg _404268_404268 ; 
   reg __404268_404268;
   reg _404269_404269 ; 
   reg __404269_404269;
   reg _404270_404270 ; 
   reg __404270_404270;
   reg _404271_404271 ; 
   reg __404271_404271;
   reg _404272_404272 ; 
   reg __404272_404272;
   reg _404273_404273 ; 
   reg __404273_404273;
   reg _404274_404274 ; 
   reg __404274_404274;
   reg _404275_404275 ; 
   reg __404275_404275;
   reg _404276_404276 ; 
   reg __404276_404276;
   reg _404277_404277 ; 
   reg __404277_404277;
   reg _404278_404278 ; 
   reg __404278_404278;
   reg _404279_404279 ; 
   reg __404279_404279;
   reg _404280_404280 ; 
   reg __404280_404280;
   reg _404281_404281 ; 
   reg __404281_404281;
   reg _404282_404282 ; 
   reg __404282_404282;
   reg _404283_404283 ; 
   reg __404283_404283;
   reg _404284_404284 ; 
   reg __404284_404284;
   reg _404285_404285 ; 
   reg __404285_404285;
   reg _404286_404286 ; 
   reg __404286_404286;
   reg _404287_404287 ; 
   reg __404287_404287;
   reg _404288_404288 ; 
   reg __404288_404288;
   reg _404289_404289 ; 
   reg __404289_404289;
   reg _404290_404290 ; 
   reg __404290_404290;
   reg _404291_404291 ; 
   reg __404291_404291;
   reg _404292_404292 ; 
   reg __404292_404292;
   reg _404293_404293 ; 
   reg __404293_404293;
   reg _404294_404294 ; 
   reg __404294_404294;
   reg _404295_404295 ; 
   reg __404295_404295;
   reg _404296_404296 ; 
   reg __404296_404296;
   reg _404297_404297 ; 
   reg __404297_404297;
   reg _404298_404298 ; 
   reg __404298_404298;
   reg _404299_404299 ; 
   reg __404299_404299;
   reg _404300_404300 ; 
   reg __404300_404300;
   reg _404301_404301 ; 
   reg __404301_404301;
   reg _404302_404302 ; 
   reg __404302_404302;
   reg _404303_404303 ; 
   reg __404303_404303;
   reg _404304_404304 ; 
   reg __404304_404304;
   reg _404305_404305 ; 
   reg __404305_404305;
   reg _404306_404306 ; 
   reg __404306_404306;
   reg _404307_404307 ; 
   reg __404307_404307;
   reg _404308_404308 ; 
   reg __404308_404308;
   reg _404309_404309 ; 
   reg __404309_404309;
   reg _404310_404310 ; 
   reg __404310_404310;
   reg _404311_404311 ; 
   reg __404311_404311;
   reg _404312_404312 ; 
   reg __404312_404312;
   reg _404313_404313 ; 
   reg __404313_404313;
   reg _404314_404314 ; 
   reg __404314_404314;
   reg _404315_404315 ; 
   reg __404315_404315;
   reg _404316_404316 ; 
   reg __404316_404316;
   reg _404317_404317 ; 
   reg __404317_404317;
   reg _404318_404318 ; 
   reg __404318_404318;
   reg _404319_404319 ; 
   reg __404319_404319;
   reg _404320_404320 ; 
   reg __404320_404320;
   reg _404321_404321 ; 
   reg __404321_404321;
   reg _404322_404322 ; 
   reg __404322_404322;
   reg _404323_404323 ; 
   reg __404323_404323;
   reg _404324_404324 ; 
   reg __404324_404324;
   reg _404325_404325 ; 
   reg __404325_404325;
   reg _404326_404326 ; 
   reg __404326_404326;
   reg _404327_404327 ; 
   reg __404327_404327;
   reg _404328_404328 ; 
   reg __404328_404328;
   reg _404329_404329 ; 
   reg __404329_404329;
   reg _404330_404330 ; 
   reg __404330_404330;
   reg _404331_404331 ; 
   reg __404331_404331;
   reg _404332_404332 ; 
   reg __404332_404332;
   reg _404333_404333 ; 
   reg __404333_404333;
   reg _404334_404334 ; 
   reg __404334_404334;
   reg _404335_404335 ; 
   reg __404335_404335;
   reg _404336_404336 ; 
   reg __404336_404336;
   reg _404337_404337 ; 
   reg __404337_404337;
   reg _404338_404338 ; 
   reg __404338_404338;
   reg _404339_404339 ; 
   reg __404339_404339;
   reg _404340_404340 ; 
   reg __404340_404340;
   reg _404341_404341 ; 
   reg __404341_404341;
   reg _404342_404342 ; 
   reg __404342_404342;
   reg _404343_404343 ; 
   reg __404343_404343;
   reg _404344_404344 ; 
   reg __404344_404344;
   reg _404345_404345 ; 
   reg __404345_404345;
   reg _404346_404346 ; 
   reg __404346_404346;
   reg _404347_404347 ; 
   reg __404347_404347;
   reg _404348_404348 ; 
   reg __404348_404348;
   reg _404349_404349 ; 
   reg __404349_404349;
   reg _404350_404350 ; 
   reg __404350_404350;
   reg _404351_404351 ; 
   reg __404351_404351;
   reg _404352_404352 ; 
   reg __404352_404352;
   reg _404353_404353 ; 
   reg __404353_404353;
   reg _404354_404354 ; 
   reg __404354_404354;
   reg _404355_404355 ; 
   reg __404355_404355;
   reg _404356_404356 ; 
   reg __404356_404356;
   reg _404357_404357 ; 
   reg __404357_404357;
   reg _404358_404358 ; 
   reg __404358_404358;
   reg _404359_404359 ; 
   reg __404359_404359;
   reg _404360_404360 ; 
   reg __404360_404360;
   reg _404361_404361 ; 
   reg __404361_404361;
   reg _404362_404362 ; 
   reg __404362_404362;
   reg _404363_404363 ; 
   reg __404363_404363;
   reg _404364_404364 ; 
   reg __404364_404364;
   reg _404365_404365 ; 
   reg __404365_404365;
   reg _404366_404366 ; 
   reg __404366_404366;
   reg _404367_404367 ; 
   reg __404367_404367;
   reg _404368_404368 ; 
   reg __404368_404368;
   reg _404369_404369 ; 
   reg __404369_404369;
   reg _404370_404370 ; 
   reg __404370_404370;
   reg _404371_404371 ; 
   reg __404371_404371;
   reg _404372_404372 ; 
   reg __404372_404372;
   reg _404373_404373 ; 
   reg __404373_404373;
   reg _404374_404374 ; 
   reg __404374_404374;
   reg _404375_404375 ; 
   reg __404375_404375;
   reg _404376_404376 ; 
   reg __404376_404376;
   reg _404377_404377 ; 
   reg __404377_404377;
   reg _404378_404378 ; 
   reg __404378_404378;
   reg _404379_404379 ; 
   reg __404379_404379;
   reg _404380_404380 ; 
   reg __404380_404380;
   reg _404381_404381 ; 
   reg __404381_404381;
   reg _404382_404382 ; 
   reg __404382_404382;
   reg _404383_404383 ; 
   reg __404383_404383;
   reg _404384_404384 ; 
   reg __404384_404384;
   reg _404385_404385 ; 
   reg __404385_404385;
   reg _404386_404386 ; 
   reg __404386_404386;
   reg _404387_404387 ; 
   reg __404387_404387;
   reg _404388_404388 ; 
   reg __404388_404388;
   reg _404389_404389 ; 
   reg __404389_404389;
   reg _404390_404390 ; 
   reg __404390_404390;
   reg _404391_404391 ; 
   reg __404391_404391;
   reg _404392_404392 ; 
   reg __404392_404392;
   reg _404393_404393 ; 
   reg __404393_404393;
   reg _404394_404394 ; 
   reg __404394_404394;
   reg _404395_404395 ; 
   reg __404395_404395;
   reg _404396_404396 ; 
   reg __404396_404396;
   reg _404397_404397 ; 
   reg __404397_404397;
   reg _404398_404398 ; 
   reg __404398_404398;
   reg _404399_404399 ; 
   reg __404399_404399;
   reg _404400_404400 ; 
   reg __404400_404400;
   reg _404401_404401 ; 
   reg __404401_404401;
   reg _404402_404402 ; 
   reg __404402_404402;
   reg _404403_404403 ; 
   reg __404403_404403;
   reg _404404_404404 ; 
   reg __404404_404404;
   reg _404405_404405 ; 
   reg __404405_404405;
   reg _404406_404406 ; 
   reg __404406_404406;
   reg _404407_404407 ; 
   reg __404407_404407;
   reg _404408_404408 ; 
   reg __404408_404408;
   reg _404409_404409 ; 
   reg __404409_404409;
   reg _404410_404410 ; 
   reg __404410_404410;
   reg _404411_404411 ; 
   reg __404411_404411;
   reg _404412_404412 ; 
   reg __404412_404412;
   reg _404413_404413 ; 
   reg __404413_404413;
   reg _404414_404414 ; 
   reg __404414_404414;
   reg _404415_404415 ; 
   reg __404415_404415;
   reg _404416_404416 ; 
   reg __404416_404416;
   reg _404417_404417 ; 
   reg __404417_404417;
   reg _404418_404418 ; 
   reg __404418_404418;
   reg _404419_404419 ; 
   reg __404419_404419;
   reg _404420_404420 ; 
   reg __404420_404420;
   reg _404421_404421 ; 
   reg __404421_404421;
   reg _404422_404422 ; 
   reg __404422_404422;
   reg _404423_404423 ; 
   reg __404423_404423;
   reg _404424_404424 ; 
   reg __404424_404424;
   reg _404425_404425 ; 
   reg __404425_404425;
   reg _404426_404426 ; 
   reg __404426_404426;
   reg _404427_404427 ; 
   reg __404427_404427;
   reg _404428_404428 ; 
   reg __404428_404428;
   reg _404429_404429 ; 
   reg __404429_404429;
   reg _404430_404430 ; 
   reg __404430_404430;
   reg _404431_404431 ; 
   reg __404431_404431;
   reg _404432_404432 ; 
   reg __404432_404432;
   reg _404433_404433 ; 
   reg __404433_404433;
   reg _404434_404434 ; 
   reg __404434_404434;
   reg _404435_404435 ; 
   reg __404435_404435;
   reg _404436_404436 ; 
   reg __404436_404436;
   reg _404437_404437 ; 
   reg __404437_404437;
   reg _404438_404438 ; 
   reg __404438_404438;
   reg _404439_404439 ; 
   reg __404439_404439;
   reg _404440_404440 ; 
   reg __404440_404440;
   reg _404441_404441 ; 
   reg __404441_404441;
   reg _404442_404442 ; 
   reg __404442_404442;
   reg _404443_404443 ; 
   reg __404443_404443;
   reg _404444_404444 ; 
   reg __404444_404444;
   reg _404445_404445 ; 
   reg __404445_404445;
   reg _404446_404446 ; 
   reg __404446_404446;
   reg _404447_404447 ; 
   reg __404447_404447;
   reg _404448_404448 ; 
   reg __404448_404448;
   reg _404449_404449 ; 
   reg __404449_404449;
   reg _404450_404450 ; 
   reg __404450_404450;
   reg _404451_404451 ; 
   reg __404451_404451;
   reg _404452_404452 ; 
   reg __404452_404452;
   reg _404453_404453 ; 
   reg __404453_404453;
   reg _404454_404454 ; 
   reg __404454_404454;
   reg _404455_404455 ; 
   reg __404455_404455;
   reg _404456_404456 ; 
   reg __404456_404456;
   reg _404457_404457 ; 
   reg __404457_404457;
   reg _404458_404458 ; 
   reg __404458_404458;
   reg _404459_404459 ; 
   reg __404459_404459;
   reg _404460_404460 ; 
   reg __404460_404460;
   reg _404461_404461 ; 
   reg __404461_404461;
   reg _404462_404462 ; 
   reg __404462_404462;
   reg _404463_404463 ; 
   reg __404463_404463;
   reg _404464_404464 ; 
   reg __404464_404464;
   reg _404465_404465 ; 
   reg __404465_404465;
   reg _404466_404466 ; 
   reg __404466_404466;
   reg _404467_404467 ; 
   reg __404467_404467;
   reg _404468_404468 ; 
   reg __404468_404468;
   reg _404469_404469 ; 
   reg __404469_404469;
   reg _404470_404470 ; 
   reg __404470_404470;
   reg _404471_404471 ; 
   reg __404471_404471;
   reg _404472_404472 ; 
   reg __404472_404472;
   reg _404473_404473 ; 
   reg __404473_404473;
   reg _404474_404474 ; 
   reg __404474_404474;
   reg _404475_404475 ; 
   reg __404475_404475;
   reg _404476_404476 ; 
   reg __404476_404476;
   reg _404477_404477 ; 
   reg __404477_404477;
   reg _404478_404478 ; 
   reg __404478_404478;
   reg _404479_404479 ; 
   reg __404479_404479;
   reg _404480_404480 ; 
   reg __404480_404480;
   reg _404481_404481 ; 
   reg __404481_404481;
   reg _404482_404482 ; 
   reg __404482_404482;
   reg _404483_404483 ; 
   reg __404483_404483;
   reg _404484_404484 ; 
   reg __404484_404484;
   reg _404485_404485 ; 
   reg __404485_404485;
   reg _404486_404486 ; 
   reg __404486_404486;
   reg _404487_404487 ; 
   reg __404487_404487;
   reg _404488_404488 ; 
   reg __404488_404488;
   reg _404489_404489 ; 
   reg __404489_404489;
   reg _404490_404490 ; 
   reg __404490_404490;
   reg _404491_404491 ; 
   reg __404491_404491;
   reg _404492_404492 ; 
   reg __404492_404492;
   reg _404493_404493 ; 
   reg __404493_404493;
   reg _404494_404494 ; 
   reg __404494_404494;
   reg _404495_404495 ; 
   reg __404495_404495;
   reg _404496_404496 ; 
   reg __404496_404496;
   reg _404497_404497 ; 
   reg __404497_404497;
   reg _404498_404498 ; 
   reg __404498_404498;
   reg _404499_404499 ; 
   reg __404499_404499;
   reg _404500_404500 ; 
   reg __404500_404500;
   reg _404501_404501 ; 
   reg __404501_404501;
   reg _404502_404502 ; 
   reg __404502_404502;
   reg _404503_404503 ; 
   reg __404503_404503;
   reg _404504_404504 ; 
   reg __404504_404504;
   reg _404505_404505 ; 
   reg __404505_404505;
   reg _404506_404506 ; 
   reg __404506_404506;
   reg _404507_404507 ; 
   reg __404507_404507;
   reg _404508_404508 ; 
   reg __404508_404508;
   reg _404509_404509 ; 
   reg __404509_404509;
   reg _404510_404510 ; 
   reg __404510_404510;
   reg _404511_404511 ; 
   reg __404511_404511;
   reg _404512_404512 ; 
   reg __404512_404512;
   reg _404513_404513 ; 
   reg __404513_404513;
   reg _404514_404514 ; 
   reg __404514_404514;
   reg _404515_404515 ; 
   reg __404515_404515;
   reg _404516_404516 ; 
   reg __404516_404516;
   reg _404517_404517 ; 
   reg __404517_404517;
   reg _404518_404518 ; 
   reg __404518_404518;
   reg _404519_404519 ; 
   reg __404519_404519;
   reg _404520_404520 ; 
   reg __404520_404520;
   reg _404521_404521 ; 
   reg __404521_404521;
   reg _404522_404522 ; 
   reg __404522_404522;
   reg _404523_404523 ; 
   reg __404523_404523;
   reg _404524_404524 ; 
   reg __404524_404524;
   reg _404525_404525 ; 
   reg __404525_404525;
   reg _404526_404526 ; 
   reg __404526_404526;
   reg _404527_404527 ; 
   reg __404527_404527;
   reg _404528_404528 ; 
   reg __404528_404528;
   reg _404529_404529 ; 
   reg __404529_404529;
   reg _404530_404530 ; 
   reg __404530_404530;
   reg _404531_404531 ; 
   reg __404531_404531;
   reg _404532_404532 ; 
   reg __404532_404532;
   reg _404533_404533 ; 
   reg __404533_404533;
   reg _404534_404534 ; 
   reg __404534_404534;
   reg _404535_404535 ; 
   reg __404535_404535;
   reg _404536_404536 ; 
   reg __404536_404536;
   reg _404537_404537 ; 
   reg __404537_404537;
   reg _404538_404538 ; 
   reg __404538_404538;
   reg _404539_404539 ; 
   reg __404539_404539;
   reg _404540_404540 ; 
   reg __404540_404540;
   reg _404541_404541 ; 
   reg __404541_404541;
   reg _404542_404542 ; 
   reg __404542_404542;
   reg _404543_404543 ; 
   reg __404543_404543;
   reg _404544_404544 ; 
   reg __404544_404544;
   reg _404545_404545 ; 
   reg __404545_404545;
   reg _404546_404546 ; 
   reg __404546_404546;
   reg _404547_404547 ; 
   reg __404547_404547;
   reg _404548_404548 ; 
   reg __404548_404548;
   reg _404549_404549 ; 
   reg __404549_404549;
   reg _404550_404550 ; 
   reg __404550_404550;
   reg _404551_404551 ; 
   reg __404551_404551;
   reg _404552_404552 ; 
   reg __404552_404552;
   reg _404553_404553 ; 
   reg __404553_404553;
   reg _404554_404554 ; 
   reg __404554_404554;
   reg _404555_404555 ; 
   reg __404555_404555;
   reg _404556_404556 ; 
   reg __404556_404556;
   reg _404557_404557 ; 
   reg __404557_404557;
   reg _404558_404558 ; 
   reg __404558_404558;
   reg _404559_404559 ; 
   reg __404559_404559;
   reg _404560_404560 ; 
   reg __404560_404560;
   reg _404561_404561 ; 
   reg __404561_404561;
   reg _404562_404562 ; 
   reg __404562_404562;
   reg _404563_404563 ; 
   reg __404563_404563;
   reg _404564_404564 ; 
   reg __404564_404564;
   reg _404565_404565 ; 
   reg __404565_404565;
   reg _404566_404566 ; 
   reg __404566_404566;
   reg _404567_404567 ; 
   reg __404567_404567;
   reg _404568_404568 ; 
   reg __404568_404568;
   reg _404569_404569 ; 
   reg __404569_404569;
   reg _404570_404570 ; 
   reg __404570_404570;
   reg _404571_404571 ; 
   reg __404571_404571;
   reg _404572_404572 ; 
   reg __404572_404572;
   reg _404573_404573 ; 
   reg __404573_404573;
   reg _404574_404574 ; 
   reg __404574_404574;
   reg _404575_404575 ; 
   reg __404575_404575;
   reg _404576_404576 ; 
   reg __404576_404576;
   reg _404577_404577 ; 
   reg __404577_404577;
   reg _404578_404578 ; 
   reg __404578_404578;
   reg _404579_404579 ; 
   reg __404579_404579;
   reg _404580_404580 ; 
   reg __404580_404580;
   reg _404581_404581 ; 
   reg __404581_404581;
   reg _404582_404582 ; 
   reg __404582_404582;
   reg _404583_404583 ; 
   reg __404583_404583;
   reg _404584_404584 ; 
   reg __404584_404584;
   reg _404585_404585 ; 
   reg __404585_404585;
   reg _404586_404586 ; 
   reg __404586_404586;
   reg _404587_404587 ; 
   reg __404587_404587;
   reg _404588_404588 ; 
   reg __404588_404588;
   reg _404589_404589 ; 
   reg __404589_404589;
   reg _404590_404590 ; 
   reg __404590_404590;
   reg _404591_404591 ; 
   reg __404591_404591;
   reg _404592_404592 ; 
   reg __404592_404592;
   reg _404593_404593 ; 
   reg __404593_404593;
   reg _404594_404594 ; 
   reg __404594_404594;
   reg _404595_404595 ; 
   reg __404595_404595;
   reg _404596_404596 ; 
   reg __404596_404596;
   reg _404597_404597 ; 
   reg __404597_404597;
   reg _404598_404598 ; 
   reg __404598_404598;
   reg _404599_404599 ; 
   reg __404599_404599;
   reg _404600_404600 ; 
   reg __404600_404600;
   reg _404601_404601 ; 
   reg __404601_404601;
   reg _404602_404602 ; 
   reg __404602_404602;
   reg _404603_404603 ; 
   reg __404603_404603;
   reg _404604_404604 ; 
   reg __404604_404604;
   reg _404605_404605 ; 
   reg __404605_404605;
   reg _404606_404606 ; 
   reg __404606_404606;
   reg _404607_404607 ; 
   reg __404607_404607;
   reg _404608_404608 ; 
   reg __404608_404608;
   reg _404609_404609 ; 
   reg __404609_404609;
   reg _404610_404610 ; 
   reg __404610_404610;
   reg _404611_404611 ; 
   reg __404611_404611;
   reg _404612_404612 ; 
   reg __404612_404612;
   reg _404613_404613 ; 
   reg __404613_404613;
   reg _404614_404614 ; 
   reg __404614_404614;
   reg _404615_404615 ; 
   reg __404615_404615;
   reg _404616_404616 ; 
   reg __404616_404616;
   reg _404617_404617 ; 
   reg __404617_404617;
   reg _404618_404618 ; 
   reg __404618_404618;
   reg _404619_404619 ; 
   reg __404619_404619;
   reg _404620_404620 ; 
   reg __404620_404620;
   reg _404621_404621 ; 
   reg __404621_404621;
   reg _404622_404622 ; 
   reg __404622_404622;
   reg _404623_404623 ; 
   reg __404623_404623;
   reg _404624_404624 ; 
   reg __404624_404624;
   reg _404625_404625 ; 
   reg __404625_404625;
   reg _404626_404626 ; 
   reg __404626_404626;
   reg _404627_404627 ; 
   reg __404627_404627;
   reg _404628_404628 ; 
   reg __404628_404628;
   reg _404629_404629 ; 
   reg __404629_404629;
   reg _404630_404630 ; 
   reg __404630_404630;
   reg _404631_404631 ; 
   reg __404631_404631;
   reg _404632_404632 ; 
   reg __404632_404632;
   reg _404633_404633 ; 
   reg __404633_404633;
   reg _404634_404634 ; 
   reg __404634_404634;
   reg _404635_404635 ; 
   reg __404635_404635;
   reg _404636_404636 ; 
   reg __404636_404636;
   reg _404637_404637 ; 
   reg __404637_404637;
   reg _404638_404638 ; 
   reg __404638_404638;
   reg _404639_404639 ; 
   reg __404639_404639;
   reg _404640_404640 ; 
   reg __404640_404640;
   reg _404641_404641 ; 
   reg __404641_404641;
   reg _404642_404642 ; 
   reg __404642_404642;
   reg _404643_404643 ; 
   reg __404643_404643;
   reg _404644_404644 ; 
   reg __404644_404644;
   reg _404645_404645 ; 
   reg __404645_404645;
   reg _404646_404646 ; 
   reg __404646_404646;
   reg _404647_404647 ; 
   reg __404647_404647;
   reg _404648_404648 ; 
   reg __404648_404648;
   reg _404649_404649 ; 
   reg __404649_404649;
   reg _404650_404650 ; 
   reg __404650_404650;
   reg _404651_404651 ; 
   reg __404651_404651;
   reg _404652_404652 ; 
   reg __404652_404652;
   reg _404653_404653 ; 
   reg __404653_404653;
   reg _404654_404654 ; 
   reg __404654_404654;
   reg _404655_404655 ; 
   reg __404655_404655;
   reg _404656_404656 ; 
   reg __404656_404656;
   reg _404657_404657 ; 
   reg __404657_404657;
   reg _404658_404658 ; 
   reg __404658_404658;
   reg _404659_404659 ; 
   reg __404659_404659;
   reg _404660_404660 ; 
   reg __404660_404660;
   reg _404661_404661 ; 
   reg __404661_404661;
   reg _404662_404662 ; 
   reg __404662_404662;
   reg _404663_404663 ; 
   reg __404663_404663;
   reg _404664_404664 ; 
   reg __404664_404664;
   reg _404665_404665 ; 
   reg __404665_404665;
   reg _404666_404666 ; 
   reg __404666_404666;
   reg _404667_404667 ; 
   reg __404667_404667;
   reg _404668_404668 ; 
   reg __404668_404668;
   reg _404669_404669 ; 
   reg __404669_404669;
   reg _404670_404670 ; 
   reg __404670_404670;
   reg _404671_404671 ; 
   reg __404671_404671;
   reg _404672_404672 ; 
   reg __404672_404672;
   reg _404673_404673 ; 
   reg __404673_404673;
   reg _404674_404674 ; 
   reg __404674_404674;
   reg _404675_404675 ; 
   reg __404675_404675;
   reg _404676_404676 ; 
   reg __404676_404676;
   reg _404677_404677 ; 
   reg __404677_404677;
   reg _404678_404678 ; 
   reg __404678_404678;
   reg _404679_404679 ; 
   reg __404679_404679;
   reg _404680_404680 ; 
   reg __404680_404680;
   reg _404681_404681 ; 
   reg __404681_404681;
   reg _404682_404682 ; 
   reg __404682_404682;
   reg _404683_404683 ; 
   reg __404683_404683;
   reg _404684_404684 ; 
   reg __404684_404684;
   reg _404685_404685 ; 
   reg __404685_404685;
   reg _404686_404686 ; 
   reg __404686_404686;
   reg _404687_404687 ; 
   reg __404687_404687;
   reg _404688_404688 ; 
   reg __404688_404688;
   reg _404689_404689 ; 
   reg __404689_404689;
   reg _404690_404690 ; 
   reg __404690_404690;
   reg _404691_404691 ; 
   reg __404691_404691;
   reg _404692_404692 ; 
   reg __404692_404692;
   reg _404693_404693 ; 
   reg __404693_404693;
   reg _404694_404694 ; 
   reg __404694_404694;
   reg _404695_404695 ; 
   reg __404695_404695;
   reg _404696_404696 ; 
   reg __404696_404696;
   reg _404697_404697 ; 
   reg __404697_404697;
   reg _404698_404698 ; 
   reg __404698_404698;
   reg _404699_404699 ; 
   reg __404699_404699;
   reg _404700_404700 ; 
   reg __404700_404700;
   reg _404701_404701 ; 
   reg __404701_404701;
   reg _404702_404702 ; 
   reg __404702_404702;
   reg _404703_404703 ; 
   reg __404703_404703;
   reg _404704_404704 ; 
   reg __404704_404704;
   reg _404705_404705 ; 
   reg __404705_404705;
   reg _404706_404706 ; 
   reg __404706_404706;
   reg _404707_404707 ; 
   reg __404707_404707;
   reg _404708_404708 ; 
   reg __404708_404708;
   reg _404709_404709 ; 
   reg __404709_404709;
   reg _404710_404710 ; 
   reg __404710_404710;
   reg _404711_404711 ; 
   reg __404711_404711;
   reg _404712_404712 ; 
   reg __404712_404712;
   reg _404713_404713 ; 
   reg __404713_404713;
   reg _404714_404714 ; 
   reg __404714_404714;
   reg _404715_404715 ; 
   reg __404715_404715;
   reg _404716_404716 ; 
   reg __404716_404716;
   reg _404717_404717 ; 
   reg __404717_404717;
   reg _404718_404718 ; 
   reg __404718_404718;
   reg _404719_404719 ; 
   reg __404719_404719;
   reg _404720_404720 ; 
   reg __404720_404720;
   reg _404721_404721 ; 
   reg __404721_404721;
   reg _404722_404722 ; 
   reg __404722_404722;
   reg _404723_404723 ; 
   reg __404723_404723;
   reg _404724_404724 ; 
   reg __404724_404724;
   reg _404725_404725 ; 
   reg __404725_404725;
   reg _404726_404726 ; 
   reg __404726_404726;
   reg _404727_404727 ; 
   reg __404727_404727;
   reg _404728_404728 ; 
   reg __404728_404728;
   reg _404729_404729 ; 
   reg __404729_404729;
   reg _404730_404730 ; 
   reg __404730_404730;
   reg _404731_404731 ; 
   reg __404731_404731;
   reg _404732_404732 ; 
   reg __404732_404732;
   reg _404733_404733 ; 
   reg __404733_404733;
   reg _404734_404734 ; 
   reg __404734_404734;
   reg _404735_404735 ; 
   reg __404735_404735;
   reg _404736_404736 ; 
   reg __404736_404736;
   reg _404737_404737 ; 
   reg __404737_404737;
   reg _404738_404738 ; 
   reg __404738_404738;
   reg _404739_404739 ; 
   reg __404739_404739;
   reg _404740_404740 ; 
   reg __404740_404740;
   reg _404741_404741 ; 
   reg __404741_404741;
   reg _404742_404742 ; 
   reg __404742_404742;
   reg _404743_404743 ; 
   reg __404743_404743;
   reg _404744_404744 ; 
   reg __404744_404744;
   reg _404745_404745 ; 
   reg __404745_404745;
   reg _404746_404746 ; 
   reg __404746_404746;
   reg _404747_404747 ; 
   reg __404747_404747;
   reg _404748_404748 ; 
   reg __404748_404748;
   reg _404749_404749 ; 
   reg __404749_404749;
   reg _404750_404750 ; 
   reg __404750_404750;
   reg _404751_404751 ; 
   reg __404751_404751;
   reg _404752_404752 ; 
   reg __404752_404752;
   reg _404753_404753 ; 
   reg __404753_404753;
   reg _404754_404754 ; 
   reg __404754_404754;
   reg _404755_404755 ; 
   reg __404755_404755;
   reg _404756_404756 ; 
   reg __404756_404756;
   reg _404757_404757 ; 
   reg __404757_404757;
   reg _404758_404758 ; 
   reg __404758_404758;
   reg _404759_404759 ; 
   reg __404759_404759;
   reg _404760_404760 ; 
   reg __404760_404760;
   reg _404761_404761 ; 
   reg __404761_404761;
   reg _404762_404762 ; 
   reg __404762_404762;
   reg _404763_404763 ; 
   reg __404763_404763;
   reg _404764_404764 ; 
   reg __404764_404764;
   reg _404765_404765 ; 
   reg __404765_404765;
   reg _404766_404766 ; 
   reg __404766_404766;
   reg _404767_404767 ; 
   reg __404767_404767;
   reg _404768_404768 ; 
   reg __404768_404768;
   reg _404769_404769 ; 
   reg __404769_404769;
   reg _404770_404770 ; 
   reg __404770_404770;
   reg _404771_404771 ; 
   reg __404771_404771;
   reg _404772_404772 ; 
   reg __404772_404772;
   reg _404773_404773 ; 
   reg __404773_404773;
   reg _404774_404774 ; 
   reg __404774_404774;
   reg _404775_404775 ; 
   reg __404775_404775;
   reg _404776_404776 ; 
   reg __404776_404776;
   reg _404777_404777 ; 
   reg __404777_404777;
   reg _404778_404778 ; 
   reg __404778_404778;
   reg _404779_404779 ; 
   reg __404779_404779;
   reg _404780_404780 ; 
   reg __404780_404780;
   reg _404781_404781 ; 
   reg __404781_404781;
   reg _404782_404782 ; 
   reg __404782_404782;
   reg _404783_404783 ; 
   reg __404783_404783;
   reg _404784_404784 ; 
   reg __404784_404784;
   reg _404785_404785 ; 
   reg __404785_404785;
   reg _404786_404786 ; 
   reg __404786_404786;
   reg _404787_404787 ; 
   reg __404787_404787;
   reg _404788_404788 ; 
   reg __404788_404788;
   reg _404789_404789 ; 
   reg __404789_404789;
   reg _404790_404790 ; 
   reg __404790_404790;
   reg _404791_404791 ; 
   reg __404791_404791;
   reg _404792_404792 ; 
   reg __404792_404792;
   reg _404793_404793 ; 
   reg __404793_404793;
   reg _404794_404794 ; 
   reg __404794_404794;
   reg _404795_404795 ; 
   reg __404795_404795;
   reg _404796_404796 ; 
   reg __404796_404796;
   reg _404797_404797 ; 
   reg __404797_404797;
   reg _404798_404798 ; 
   reg __404798_404798;
   reg _404799_404799 ; 
   reg __404799_404799;
   reg _404800_404800 ; 
   reg __404800_404800;
   reg _404801_404801 ; 
   reg __404801_404801;
   reg _404802_404802 ; 
   reg __404802_404802;
   reg _404803_404803 ; 
   reg __404803_404803;
   reg _404804_404804 ; 
   reg __404804_404804;
   reg _404805_404805 ; 
   reg __404805_404805;
   reg _404806_404806 ; 
   reg __404806_404806;
   reg _404807_404807 ; 
   reg __404807_404807;
   reg _404808_404808 ; 
   reg __404808_404808;
   reg _404809_404809 ; 
   reg __404809_404809;
   reg _404810_404810 ; 
   reg __404810_404810;
   reg _404811_404811 ; 
   reg __404811_404811;
   reg _404812_404812 ; 
   reg __404812_404812;
   reg _404813_404813 ; 
   reg __404813_404813;
   reg _404814_404814 ; 
   reg __404814_404814;
   reg _404815_404815 ; 
   reg __404815_404815;
   reg _404816_404816 ; 
   reg __404816_404816;
   reg _404817_404817 ; 
   reg __404817_404817;
   reg _404818_404818 ; 
   reg __404818_404818;
   reg _404819_404819 ; 
   reg __404819_404819;
   reg _404820_404820 ; 
   reg __404820_404820;
   reg _404821_404821 ; 
   reg __404821_404821;
   reg _404822_404822 ; 
   reg __404822_404822;
   reg _404823_404823 ; 
   reg __404823_404823;
   reg _404824_404824 ; 
   reg __404824_404824;
   reg _404825_404825 ; 
   reg __404825_404825;
   reg _404826_404826 ; 
   reg __404826_404826;
   reg _404827_404827 ; 
   reg __404827_404827;
   reg _404828_404828 ; 
   reg __404828_404828;
   reg _404829_404829 ; 
   reg __404829_404829;
   reg _404830_404830 ; 
   reg __404830_404830;
   reg _404831_404831 ; 
   reg __404831_404831;
   reg _404832_404832 ; 
   reg __404832_404832;
   reg _404833_404833 ; 
   reg __404833_404833;
   reg _404834_404834 ; 
   reg __404834_404834;
   reg _404835_404835 ; 
   reg __404835_404835;
   reg _404836_404836 ; 
   reg __404836_404836;
   reg _404837_404837 ; 
   reg __404837_404837;
   reg _404838_404838 ; 
   reg __404838_404838;
   reg _404839_404839 ; 
   reg __404839_404839;
   reg _404840_404840 ; 
   reg __404840_404840;
   reg _404841_404841 ; 
   reg __404841_404841;
   reg _404842_404842 ; 
   reg __404842_404842;
   reg _404843_404843 ; 
   reg __404843_404843;
   reg _404844_404844 ; 
   reg __404844_404844;
   reg _404845_404845 ; 
   reg __404845_404845;
   reg _404846_404846 ; 
   reg __404846_404846;
   reg _404847_404847 ; 
   reg __404847_404847;
   reg _404848_404848 ; 
   reg __404848_404848;
   reg _404849_404849 ; 
   reg __404849_404849;
   reg _404850_404850 ; 
   reg __404850_404850;
   reg _404851_404851 ; 
   reg __404851_404851;
   reg _404852_404852 ; 
   reg __404852_404852;
   reg _404853_404853 ; 
   reg __404853_404853;
   reg _404854_404854 ; 
   reg __404854_404854;
   reg _404855_404855 ; 
   reg __404855_404855;
   reg _404856_404856 ; 
   reg __404856_404856;
   reg _404857_404857 ; 
   reg __404857_404857;
   reg _404858_404858 ; 
   reg __404858_404858;
   reg _404859_404859 ; 
   reg __404859_404859;
   reg _404860_404860 ; 
   reg __404860_404860;
   reg _404861_404861 ; 
   reg __404861_404861;
   reg _404862_404862 ; 
   reg __404862_404862;
   reg _404863_404863 ; 
   reg __404863_404863;
   reg _404864_404864 ; 
   reg __404864_404864;
   reg _404865_404865 ; 
   reg __404865_404865;
   reg _404866_404866 ; 
   reg __404866_404866;
   reg _404867_404867 ; 
   reg __404867_404867;
   reg _404868_404868 ; 
   reg __404868_404868;
   reg _404869_404869 ; 
   reg __404869_404869;
   reg _404870_404870 ; 
   reg __404870_404870;
   reg _404871_404871 ; 
   reg __404871_404871;
   reg _404872_404872 ; 
   reg __404872_404872;
   reg _404873_404873 ; 
   reg __404873_404873;
   reg _404874_404874 ; 
   reg __404874_404874;
   reg _404875_404875 ; 
   reg __404875_404875;
   reg _404876_404876 ; 
   reg __404876_404876;
   reg _404877_404877 ; 
   reg __404877_404877;
   reg _404878_404878 ; 
   reg __404878_404878;
   reg _404879_404879 ; 
   reg __404879_404879;
   reg _404880_404880 ; 
   reg __404880_404880;
   reg _404881_404881 ; 
   reg __404881_404881;
   reg _404882_404882 ; 
   reg __404882_404882;
   reg _404883_404883 ; 
   reg __404883_404883;
   reg _404884_404884 ; 
   reg __404884_404884;
   reg _404885_404885 ; 
   reg __404885_404885;
   reg _404886_404886 ; 
   reg __404886_404886;
   reg _404887_404887 ; 
   reg __404887_404887;
   reg _404888_404888 ; 
   reg __404888_404888;
   reg _404889_404889 ; 
   reg __404889_404889;
   reg _404890_404890 ; 
   reg __404890_404890;
   reg _404891_404891 ; 
   reg __404891_404891;
   reg _404892_404892 ; 
   reg __404892_404892;
   reg _404893_404893 ; 
   reg __404893_404893;
   reg _404894_404894 ; 
   reg __404894_404894;
   reg _404895_404895 ; 
   reg __404895_404895;
   reg _404896_404896 ; 
   reg __404896_404896;
   reg _404897_404897 ; 
   reg __404897_404897;
   reg _404898_404898 ; 
   reg __404898_404898;
   reg _404899_404899 ; 
   reg __404899_404899;
   reg _404900_404900 ; 
   reg __404900_404900;
   reg _404901_404901 ; 
   reg __404901_404901;
   reg _404902_404902 ; 
   reg __404902_404902;
   reg _404903_404903 ; 
   reg __404903_404903;
   reg _404904_404904 ; 
   reg __404904_404904;
   reg _404905_404905 ; 
   reg __404905_404905;
   reg _404906_404906 ; 
   reg __404906_404906;
   reg _404907_404907 ; 
   reg __404907_404907;
   reg _404908_404908 ; 
   reg __404908_404908;
   reg _404909_404909 ; 
   reg __404909_404909;
   reg _404910_404910 ; 
   reg __404910_404910;
   reg _404911_404911 ; 
   reg __404911_404911;
   reg _404912_404912 ; 
   reg __404912_404912;
   reg _404913_404913 ; 
   reg __404913_404913;
   reg _404914_404914 ; 
   reg __404914_404914;
   reg _404915_404915 ; 
   reg __404915_404915;
   reg _404916_404916 ; 
   reg __404916_404916;
   reg _404917_404917 ; 
   reg __404917_404917;
   reg _404918_404918 ; 
   reg __404918_404918;
   reg _404919_404919 ; 
   reg __404919_404919;
   reg _404920_404920 ; 
   reg __404920_404920;
   reg _404921_404921 ; 
   reg __404921_404921;
   reg _404922_404922 ; 
   reg __404922_404922;
   reg _404923_404923 ; 
   reg __404923_404923;
   reg _404924_404924 ; 
   reg __404924_404924;
   reg _404925_404925 ; 
   reg __404925_404925;
   reg _404926_404926 ; 
   reg __404926_404926;
   reg _404927_404927 ; 
   reg __404927_404927;
   reg _404928_404928 ; 
   reg __404928_404928;
   reg _404929_404929 ; 
   reg __404929_404929;
   reg _404930_404930 ; 
   reg __404930_404930;
   reg _404931_404931 ; 
   reg __404931_404931;
   reg _404932_404932 ; 
   reg __404932_404932;
   reg _404933_404933 ; 
   reg __404933_404933;
   reg _404934_404934 ; 
   reg __404934_404934;
   reg _404935_404935 ; 
   reg __404935_404935;
   reg _404936_404936 ; 
   reg __404936_404936;
   reg _404937_404937 ; 
   reg __404937_404937;
   reg _404938_404938 ; 
   reg __404938_404938;
   reg _404939_404939 ; 
   reg __404939_404939;
   reg _404940_404940 ; 
   reg __404940_404940;
   reg _404941_404941 ; 
   reg __404941_404941;
   reg _404942_404942 ; 
   reg __404942_404942;
   reg _404943_404943 ; 
   reg __404943_404943;
   reg _404944_404944 ; 
   reg __404944_404944;
   reg _404945_404945 ; 
   reg __404945_404945;
   reg _404946_404946 ; 
   reg __404946_404946;
   reg _404947_404947 ; 
   reg __404947_404947;
   reg _404948_404948 ; 
   reg __404948_404948;
   reg _404949_404949 ; 
   reg __404949_404949;
   reg _404950_404950 ; 
   reg __404950_404950;
   reg _404951_404951 ; 
   reg __404951_404951;
   reg _404952_404952 ; 
   reg __404952_404952;
   reg _404953_404953 ; 
   reg __404953_404953;
   reg _404954_404954 ; 
   reg __404954_404954;
   reg _404955_404955 ; 
   reg __404955_404955;
   reg _404956_404956 ; 
   reg __404956_404956;
   reg _404957_404957 ; 
   reg __404957_404957;
   reg _404958_404958 ; 
   reg __404958_404958;
   reg _404959_404959 ; 
   reg __404959_404959;
   reg _404960_404960 ; 
   reg __404960_404960;
   reg _404961_404961 ; 
   reg __404961_404961;
   reg _404962_404962 ; 
   reg __404962_404962;
   reg _404963_404963 ; 
   reg __404963_404963;
   reg _404964_404964 ; 
   reg __404964_404964;
   reg _404965_404965 ; 
   reg __404965_404965;
   reg _404966_404966 ; 
   reg __404966_404966;
   reg _404967_404967 ; 
   reg __404967_404967;
   reg _404968_404968 ; 
   reg __404968_404968;
   reg _404969_404969 ; 
   reg __404969_404969;
   reg _404970_404970 ; 
   reg __404970_404970;
   reg _404971_404971 ; 
   reg __404971_404971;
   reg _404972_404972 ; 
   reg __404972_404972;
   reg _404973_404973 ; 
   reg __404973_404973;
   reg _404974_404974 ; 
   reg __404974_404974;
   reg _404975_404975 ; 
   reg __404975_404975;
   reg _404976_404976 ; 
   reg __404976_404976;
   reg _404977_404977 ; 
   reg __404977_404977;
   reg _404978_404978 ; 
   reg __404978_404978;
   reg _404979_404979 ; 
   reg __404979_404979;
   reg _404980_404980 ; 
   reg __404980_404980;
   reg _404981_404981 ; 
   reg __404981_404981;
   reg _404982_404982 ; 
   reg __404982_404982;
   reg _404983_404983 ; 
   reg __404983_404983;
   reg _404984_404984 ; 
   reg __404984_404984;
   reg _404985_404985 ; 
   reg __404985_404985;
   reg _404986_404986 ; 
   reg __404986_404986;
   reg _404987_404987 ; 
   reg __404987_404987;
   reg _404988_404988 ; 
   reg __404988_404988;
   reg _404989_404989 ; 
   reg __404989_404989;
   reg _404990_404990 ; 
   reg __404990_404990;
   reg _404991_404991 ; 
   reg __404991_404991;
   reg _404992_404992 ; 
   reg __404992_404992;
   reg _404993_404993 ; 
   reg __404993_404993;
   reg _404994_404994 ; 
   reg __404994_404994;
   reg _404995_404995 ; 
   reg __404995_404995;
   reg _404996_404996 ; 
   reg __404996_404996;
   reg _404997_404997 ; 
   reg __404997_404997;
   reg _404998_404998 ; 
   reg __404998_404998;
   reg _404999_404999 ; 
   reg __404999_404999;
   reg _405000_405000 ; 
   reg __405000_405000;
   reg _405001_405001 ; 
   reg __405001_405001;
   reg _405002_405002 ; 
   reg __405002_405002;
   reg _405003_405003 ; 
   reg __405003_405003;
   reg _405004_405004 ; 
   reg __405004_405004;
   reg _405005_405005 ; 
   reg __405005_405005;
   reg _405006_405006 ; 
   reg __405006_405006;
   reg _405007_405007 ; 
   reg __405007_405007;
   reg _405008_405008 ; 
   reg __405008_405008;
   reg _405009_405009 ; 
   reg __405009_405009;
   reg _405010_405010 ; 
   reg __405010_405010;
   reg _405011_405011 ; 
   reg __405011_405011;
   reg _405012_405012 ; 
   reg __405012_405012;
   reg _405013_405013 ; 
   reg __405013_405013;
   reg _405014_405014 ; 
   reg __405014_405014;
   reg _405015_405015 ; 
   reg __405015_405015;
   reg _405016_405016 ; 
   reg __405016_405016;
   reg _405017_405017 ; 
   reg __405017_405017;
   reg _405018_405018 ; 
   reg __405018_405018;
   reg _405019_405019 ; 
   reg __405019_405019;
   reg _405020_405020 ; 
   reg __405020_405020;
   reg _405021_405021 ; 
   reg __405021_405021;
   reg _405022_405022 ; 
   reg __405022_405022;
   reg _405023_405023 ; 
   reg __405023_405023;
   reg _405024_405024 ; 
   reg __405024_405024;
   reg _405025_405025 ; 
   reg __405025_405025;
   reg _405026_405026 ; 
   reg __405026_405026;
   reg _405027_405027 ; 
   reg __405027_405027;
   reg _405028_405028 ; 
   reg __405028_405028;
   reg _405029_405029 ; 
   reg __405029_405029;
   reg _405030_405030 ; 
   reg __405030_405030;
   reg _405031_405031 ; 
   reg __405031_405031;
   reg _405032_405032 ; 
   reg __405032_405032;
   reg _405033_405033 ; 
   reg __405033_405033;
   reg _405034_405034 ; 
   reg __405034_405034;
   reg _405035_405035 ; 
   reg __405035_405035;
   reg _405036_405036 ; 
   reg __405036_405036;
   reg _405037_405037 ; 
   reg __405037_405037;
   reg _405038_405038 ; 
   reg __405038_405038;
   reg _405039_405039 ; 
   reg __405039_405039;
   reg _405040_405040 ; 
   reg __405040_405040;
   reg _405041_405041 ; 
   reg __405041_405041;
   reg _405042_405042 ; 
   reg __405042_405042;
   reg _405043_405043 ; 
   reg __405043_405043;
   reg _405044_405044 ; 
   reg __405044_405044;
   reg _405045_405045 ; 
   reg __405045_405045;
   reg _405046_405046 ; 
   reg __405046_405046;
   reg _405047_405047 ; 
   reg __405047_405047;
   reg _405048_405048 ; 
   reg __405048_405048;
   reg _405049_405049 ; 
   reg __405049_405049;
   reg _405050_405050 ; 
   reg __405050_405050;
   reg _405051_405051 ; 
   reg __405051_405051;
   reg _405052_405052 ; 
   reg __405052_405052;
   reg _405053_405053 ; 
   reg __405053_405053;
   reg _405054_405054 ; 
   reg __405054_405054;
   reg _405055_405055 ; 
   reg __405055_405055;
   reg _405056_405056 ; 
   reg __405056_405056;
   reg _405057_405057 ; 
   reg __405057_405057;
   reg _405058_405058 ; 
   reg __405058_405058;
   reg _405059_405059 ; 
   reg __405059_405059;
   reg _405060_405060 ; 
   reg __405060_405060;
   reg _405061_405061 ; 
   reg __405061_405061;
   reg _405062_405062 ; 
   reg __405062_405062;
   reg _405063_405063 ; 
   reg __405063_405063;
   reg _405064_405064 ; 
   reg __405064_405064;
   reg _405065_405065 ; 
   reg __405065_405065;
   reg _405066_405066 ; 
   reg __405066_405066;
   reg _405067_405067 ; 
   reg __405067_405067;
   reg _405068_405068 ; 
   reg __405068_405068;
   reg _405069_405069 ; 
   reg __405069_405069;
   reg _405070_405070 ; 
   reg __405070_405070;
   reg _405071_405071 ; 
   reg __405071_405071;
   reg _405072_405072 ; 
   reg __405072_405072;
   reg _405073_405073 ; 
   reg __405073_405073;
   reg _405074_405074 ; 
   reg __405074_405074;
   reg _405075_405075 ; 
   reg __405075_405075;
   reg _405076_405076 ; 
   reg __405076_405076;
   reg _405077_405077 ; 
   reg __405077_405077;
   reg _405078_405078 ; 
   reg __405078_405078;
   reg _405079_405079 ; 
   reg __405079_405079;
   reg _405080_405080 ; 
   reg __405080_405080;
   reg _405081_405081 ; 
   reg __405081_405081;
   reg _405082_405082 ; 
   reg __405082_405082;
   reg _405083_405083 ; 
   reg __405083_405083;
   reg _405084_405084 ; 
   reg __405084_405084;
   reg _405085_405085 ; 
   reg __405085_405085;
   reg _405086_405086 ; 
   reg __405086_405086;
   reg _405087_405087 ; 
   reg __405087_405087;
   reg _405088_405088 ; 
   reg __405088_405088;
   reg _405089_405089 ; 
   reg __405089_405089;
   reg _405090_405090 ; 
   reg __405090_405090;
   reg _405091_405091 ; 
   reg __405091_405091;
   reg _405092_405092 ; 
   reg __405092_405092;
   reg _405093_405093 ; 
   reg __405093_405093;
   reg _405094_405094 ; 
   reg __405094_405094;
   reg _405095_405095 ; 
   reg __405095_405095;
   reg _405096_405096 ; 
   reg __405096_405096;
   reg _405097_405097 ; 
   reg __405097_405097;
   reg _405098_405098 ; 
   reg __405098_405098;
   reg _405099_405099 ; 
   reg __405099_405099;
   reg _405100_405100 ; 
   reg __405100_405100;
   reg _405101_405101 ; 
   reg __405101_405101;
   reg _405102_405102 ; 
   reg __405102_405102;
   reg _405103_405103 ; 
   reg __405103_405103;
   reg _405104_405104 ; 
   reg __405104_405104;
   reg _405105_405105 ; 
   reg __405105_405105;
   reg _405106_405106 ; 
   reg __405106_405106;
   reg _405107_405107 ; 
   reg __405107_405107;
   reg _405108_405108 ; 
   reg __405108_405108;
   reg _405109_405109 ; 
   reg __405109_405109;
   reg _405110_405110 ; 
   reg __405110_405110;
   reg _405111_405111 ; 
   reg __405111_405111;
   reg _405112_405112 ; 
   reg __405112_405112;
   reg _405113_405113 ; 
   reg __405113_405113;
   reg _405114_405114 ; 
   reg __405114_405114;
   reg _405115_405115 ; 
   reg __405115_405115;
   reg _405116_405116 ; 
   reg __405116_405116;
   reg _405117_405117 ; 
   reg __405117_405117;
   reg _405118_405118 ; 
   reg __405118_405118;
   reg _405119_405119 ; 
   reg __405119_405119;
   reg _405120_405120 ; 
   reg __405120_405120;
   reg _405121_405121 ; 
   reg __405121_405121;
   reg _405122_405122 ; 
   reg __405122_405122;
   reg _405123_405123 ; 
   reg __405123_405123;
   reg _405124_405124 ; 
   reg __405124_405124;
   reg _405125_405125 ; 
   reg __405125_405125;
   reg _405126_405126 ; 
   reg __405126_405126;
   reg _405127_405127 ; 
   reg __405127_405127;
   reg _405128_405128 ; 
   reg __405128_405128;
   reg _405129_405129 ; 
   reg __405129_405129;
   reg _405130_405130 ; 
   reg __405130_405130;
   reg _405131_405131 ; 
   reg __405131_405131;
   reg _405132_405132 ; 
   reg __405132_405132;
   reg _405133_405133 ; 
   reg __405133_405133;
   reg _405134_405134 ; 
   reg __405134_405134;
   reg _405135_405135 ; 
   reg __405135_405135;
   reg _405136_405136 ; 
   reg __405136_405136;
   reg _405137_405137 ; 
   reg __405137_405137;
   reg _405138_405138 ; 
   reg __405138_405138;
   reg _405139_405139 ; 
   reg __405139_405139;
   reg _405140_405140 ; 
   reg __405140_405140;
   reg _405141_405141 ; 
   reg __405141_405141;
   reg _405142_405142 ; 
   reg __405142_405142;
   reg _405143_405143 ; 
   reg __405143_405143;
   reg _405144_405144 ; 
   reg __405144_405144;
   reg _405145_405145 ; 
   reg __405145_405145;
   reg _405146_405146 ; 
   reg __405146_405146;
   reg _405147_405147 ; 
   reg __405147_405147;
   reg _405148_405148 ; 
   reg __405148_405148;
   reg _405149_405149 ; 
   reg __405149_405149;
   reg _405150_405150 ; 
   reg __405150_405150;
   reg _405151_405151 ; 
   reg __405151_405151;
   reg _405152_405152 ; 
   reg __405152_405152;
   reg _405153_405153 ; 
   reg __405153_405153;
   reg _405154_405154 ; 
   reg __405154_405154;
   reg _405155_405155 ; 
   reg __405155_405155;
   reg _405156_405156 ; 
   reg __405156_405156;
   reg _405157_405157 ; 
   reg __405157_405157;
   reg _405158_405158 ; 
   reg __405158_405158;
   reg _405159_405159 ; 
   reg __405159_405159;
   reg _405160_405160 ; 
   reg __405160_405160;
   reg _405161_405161 ; 
   reg __405161_405161;
   reg _405162_405162 ; 
   reg __405162_405162;
   reg _405163_405163 ; 
   reg __405163_405163;
   reg _405164_405164 ; 
   reg __405164_405164;
   reg _405165_405165 ; 
   reg __405165_405165;
   reg _405166_405166 ; 
   reg __405166_405166;
   reg _405167_405167 ; 
   reg __405167_405167;
   reg _405168_405168 ; 
   reg __405168_405168;
   reg _405169_405169 ; 
   reg __405169_405169;
   reg _405170_405170 ; 
   reg __405170_405170;
   reg _405171_405171 ; 
   reg __405171_405171;
   reg _405172_405172 ; 
   reg __405172_405172;
   reg _405173_405173 ; 
   reg __405173_405173;
   reg _405174_405174 ; 
   reg __405174_405174;
   reg _405175_405175 ; 
   reg __405175_405175;
   reg _405176_405176 ; 
   reg __405176_405176;
   reg _405177_405177 ; 
   reg __405177_405177;
   reg _405178_405178 ; 
   reg __405178_405178;
   reg _405179_405179 ; 
   reg __405179_405179;
   reg _405180_405180 ; 
   reg __405180_405180;
   reg _405181_405181 ; 
   reg __405181_405181;
   reg _405182_405182 ; 
   reg __405182_405182;
   reg _405183_405183 ; 
   reg __405183_405183;
   reg _405184_405184 ; 
   reg __405184_405184;
   reg _405185_405185 ; 
   reg __405185_405185;
   reg _405186_405186 ; 
   reg __405186_405186;
   reg _405187_405187 ; 
   reg __405187_405187;
   reg _405188_405188 ; 
   reg __405188_405188;
   reg _405189_405189 ; 
   reg __405189_405189;
   reg _405190_405190 ; 
   reg __405190_405190;
   reg _405191_405191 ; 
   reg __405191_405191;
   reg _405192_405192 ; 
   reg __405192_405192;
   reg _405193_405193 ; 
   reg __405193_405193;
   reg _405194_405194 ; 
   reg __405194_405194;
   reg _405195_405195 ; 
   reg __405195_405195;
   reg _405196_405196 ; 
   reg __405196_405196;
   reg _405197_405197 ; 
   reg __405197_405197;
   reg _405198_405198 ; 
   reg __405198_405198;
   reg _405199_405199 ; 
   reg __405199_405199;
   reg _405200_405200 ; 
   reg __405200_405200;
   reg _405201_405201 ; 
   reg __405201_405201;
   reg _405202_405202 ; 
   reg __405202_405202;
   reg _405203_405203 ; 
   reg __405203_405203;
   reg _405204_405204 ; 
   reg __405204_405204;
   reg _405205_405205 ; 
   reg __405205_405205;
   reg _405206_405206 ; 
   reg __405206_405206;
   reg _405207_405207 ; 
   reg __405207_405207;
   reg _405208_405208 ; 
   reg __405208_405208;
   reg _405209_405209 ; 
   reg __405209_405209;
   reg _405210_405210 ; 
   reg __405210_405210;
   reg _405211_405211 ; 
   reg __405211_405211;
   reg _405212_405212 ; 
   reg __405212_405212;
   reg _405213_405213 ; 
   reg __405213_405213;
   reg _405214_405214 ; 
   reg __405214_405214;
   reg _405215_405215 ; 
   reg __405215_405215;
   reg _405216_405216 ; 
   reg __405216_405216;
   reg _405217_405217 ; 
   reg __405217_405217;
   reg _405218_405218 ; 
   reg __405218_405218;
   reg _405219_405219 ; 
   reg __405219_405219;
   reg _405220_405220 ; 
   reg __405220_405220;
   reg _405221_405221 ; 
   reg __405221_405221;
   reg _405222_405222 ; 
   reg __405222_405222;
   reg _405223_405223 ; 
   reg __405223_405223;
   reg _405224_405224 ; 
   reg __405224_405224;
   reg _405225_405225 ; 
   reg __405225_405225;
   reg _405226_405226 ; 
   reg __405226_405226;
   reg _405227_405227 ; 
   reg __405227_405227;
   reg _405228_405228 ; 
   reg __405228_405228;
   reg _405229_405229 ; 
   reg __405229_405229;
   reg _405230_405230 ; 
   reg __405230_405230;
   reg _405231_405231 ; 
   reg __405231_405231;
   reg _405232_405232 ; 
   reg __405232_405232;
   reg _405233_405233 ; 
   reg __405233_405233;
   reg _405234_405234 ; 
   reg __405234_405234;
   reg _405235_405235 ; 
   reg __405235_405235;
   reg _405236_405236 ; 
   reg __405236_405236;
   reg _405237_405237 ; 
   reg __405237_405237;
   reg _405238_405238 ; 
   reg __405238_405238;
   reg _405239_405239 ; 
   reg __405239_405239;
   reg _405240_405240 ; 
   reg __405240_405240;
   reg _405241_405241 ; 
   reg __405241_405241;
   reg _405242_405242 ; 
   reg __405242_405242;
   reg _405243_405243 ; 
   reg __405243_405243;
   reg _405244_405244 ; 
   reg __405244_405244;
   reg _405245_405245 ; 
   reg __405245_405245;
   reg _405246_405246 ; 
   reg __405246_405246;
   reg _405247_405247 ; 
   reg __405247_405247;
   reg _405248_405248 ; 
   reg __405248_405248;
   reg _405249_405249 ; 
   reg __405249_405249;
   reg _405250_405250 ; 
   reg __405250_405250;
   reg _405251_405251 ; 
   reg __405251_405251;
   reg _405252_405252 ; 
   reg __405252_405252;
   reg _405253_405253 ; 
   reg __405253_405253;
   reg _405254_405254 ; 
   reg __405254_405254;
   reg _405255_405255 ; 
   reg __405255_405255;
   reg _405256_405256 ; 
   reg __405256_405256;
   reg _405257_405257 ; 
   reg __405257_405257;
   reg _405258_405258 ; 
   reg __405258_405258;
   reg _405259_405259 ; 
   reg __405259_405259;
   reg _405260_405260 ; 
   reg __405260_405260;
   reg _405261_405261 ; 
   reg __405261_405261;
   reg _405262_405262 ; 
   reg __405262_405262;
   reg _405263_405263 ; 
   reg __405263_405263;
   reg _405264_405264 ; 
   reg __405264_405264;
   reg _405265_405265 ; 
   reg __405265_405265;
   reg _405266_405266 ; 
   reg __405266_405266;
   reg _405267_405267 ; 
   reg __405267_405267;
   reg _405268_405268 ; 
   reg __405268_405268;
   reg _405269_405269 ; 
   reg __405269_405269;
   reg _405270_405270 ; 
   reg __405270_405270;
   reg _405271_405271 ; 
   reg __405271_405271;
   reg _405272_405272 ; 
   reg __405272_405272;
   reg _405273_405273 ; 
   reg __405273_405273;
   reg _405274_405274 ; 
   reg __405274_405274;
   reg _405275_405275 ; 
   reg __405275_405275;
   reg _405276_405276 ; 
   reg __405276_405276;
   reg _405277_405277 ; 
   reg __405277_405277;
   reg _405278_405278 ; 
   reg __405278_405278;
   reg _405279_405279 ; 
   reg __405279_405279;
   reg _405280_405280 ; 
   reg __405280_405280;
   reg _405281_405281 ; 
   reg __405281_405281;
   reg _405282_405282 ; 
   reg __405282_405282;
   reg _405283_405283 ; 
   reg __405283_405283;
   reg _405284_405284 ; 
   reg __405284_405284;
   reg _405285_405285 ; 
   reg __405285_405285;
   reg _405286_405286 ; 
   reg __405286_405286;
   reg _405287_405287 ; 
   reg __405287_405287;
   reg _405288_405288 ; 
   reg __405288_405288;
   reg _405289_405289 ; 
   reg __405289_405289;
   reg _405290_405290 ; 
   reg __405290_405290;
   reg _405291_405291 ; 
   reg __405291_405291;
   reg _405292_405292 ; 
   reg __405292_405292;
   reg _405293_405293 ; 
   reg __405293_405293;
   reg _405294_405294 ; 
   reg __405294_405294;
   reg _405295_405295 ; 
   reg __405295_405295;
   reg _405296_405296 ; 
   reg __405296_405296;
   reg _405297_405297 ; 
   reg __405297_405297;
   reg _405298_405298 ; 
   reg __405298_405298;
   reg _405299_405299 ; 
   reg __405299_405299;
   reg _405300_405300 ; 
   reg __405300_405300;
   reg _405301_405301 ; 
   reg __405301_405301;
   reg _405302_405302 ; 
   reg __405302_405302;
   reg _405303_405303 ; 
   reg __405303_405303;
   reg _405304_405304 ; 
   reg __405304_405304;
   reg _405305_405305 ; 
   reg __405305_405305;
   reg _405306_405306 ; 
   reg __405306_405306;
   reg _405307_405307 ; 
   reg __405307_405307;
   reg _405308_405308 ; 
   reg __405308_405308;
   reg _405309_405309 ; 
   reg __405309_405309;
   reg _405310_405310 ; 
   reg __405310_405310;
   reg _405311_405311 ; 
   reg __405311_405311;
   reg _405312_405312 ; 
   reg __405312_405312;
   reg _405313_405313 ; 
   reg __405313_405313;
   reg _405314_405314 ; 
   reg __405314_405314;
   reg _405315_405315 ; 
   reg __405315_405315;
   reg _405316_405316 ; 
   reg __405316_405316;
   reg _405317_405317 ; 
   reg __405317_405317;
   reg _405318_405318 ; 
   reg __405318_405318;
   reg _405319_405319 ; 
   reg __405319_405319;
   reg _405320_405320 ; 
   reg __405320_405320;
   reg _405321_405321 ; 
   reg __405321_405321;
   reg _405322_405322 ; 
   reg __405322_405322;
   reg _405323_405323 ; 
   reg __405323_405323;
   reg _405324_405324 ; 
   reg __405324_405324;
   reg _405325_405325 ; 
   reg __405325_405325;
   reg _405326_405326 ; 
   reg __405326_405326;
   reg _405327_405327 ; 
   reg __405327_405327;
   reg _405328_405328 ; 
   reg __405328_405328;
   reg _405329_405329 ; 
   reg __405329_405329;
   reg _405330_405330 ; 
   reg __405330_405330;
   reg _405331_405331 ; 
   reg __405331_405331;
   reg _405332_405332 ; 
   reg __405332_405332;
   reg _405333_405333 ; 
   reg __405333_405333;
   reg _405334_405334 ; 
   reg __405334_405334;
   reg _405335_405335 ; 
   reg __405335_405335;
   reg _405336_405336 ; 
   reg __405336_405336;
   reg _405337_405337 ; 
   reg __405337_405337;
   reg _405338_405338 ; 
   reg __405338_405338;
   reg _405339_405339 ; 
   reg __405339_405339;
   reg _405340_405340 ; 
   reg __405340_405340;
   reg _405341_405341 ; 
   reg __405341_405341;
   reg _405342_405342 ; 
   reg __405342_405342;
   reg _405343_405343 ; 
   reg __405343_405343;
   reg _405344_405344 ; 
   reg __405344_405344;
   reg _405345_405345 ; 
   reg __405345_405345;
   reg _405346_405346 ; 
   reg __405346_405346;
   reg _405347_405347 ; 
   reg __405347_405347;
   reg _405348_405348 ; 
   reg __405348_405348;
   reg _405349_405349 ; 
   reg __405349_405349;
   reg _405350_405350 ; 
   reg __405350_405350;
   reg _405351_405351 ; 
   reg __405351_405351;
   reg _405352_405352 ; 
   reg __405352_405352;
   reg _405353_405353 ; 
   reg __405353_405353;
   reg _405354_405354 ; 
   reg __405354_405354;
   reg _405355_405355 ; 
   reg __405355_405355;
   reg _405356_405356 ; 
   reg __405356_405356;
   reg _405357_405357 ; 
   reg __405357_405357;
   reg _405358_405358 ; 
   reg __405358_405358;
   reg _405359_405359 ; 
   reg __405359_405359;
   reg _405360_405360 ; 
   reg __405360_405360;
   reg _405361_405361 ; 
   reg __405361_405361;
   reg _405362_405362 ; 
   reg __405362_405362;
   reg _405363_405363 ; 
   reg __405363_405363;
   reg _405364_405364 ; 
   reg __405364_405364;
   reg _405365_405365 ; 
   reg __405365_405365;
   reg _405366_405366 ; 
   reg __405366_405366;
   reg _405367_405367 ; 
   reg __405367_405367;
   reg _405368_405368 ; 
   reg __405368_405368;
   reg _405369_405369 ; 
   reg __405369_405369;
   reg _405370_405370 ; 
   reg __405370_405370;
   reg _405371_405371 ; 
   reg __405371_405371;
   reg _405372_405372 ; 
   reg __405372_405372;
   reg _405373_405373 ; 
   reg __405373_405373;
   reg _405374_405374 ; 
   reg __405374_405374;
   reg _405375_405375 ; 
   reg __405375_405375;
   reg _405376_405376 ; 
   reg __405376_405376;
   reg _405377_405377 ; 
   reg __405377_405377;
   reg _405378_405378 ; 
   reg __405378_405378;
   reg _405379_405379 ; 
   reg __405379_405379;
   reg _405380_405380 ; 
   reg __405380_405380;
   reg _405381_405381 ; 
   reg __405381_405381;
   reg _405382_405382 ; 
   reg __405382_405382;
   reg _405383_405383 ; 
   reg __405383_405383;
   reg _405384_405384 ; 
   reg __405384_405384;
   reg _405385_405385 ; 
   reg __405385_405385;
   reg _405386_405386 ; 
   reg __405386_405386;
   reg _405387_405387 ; 
   reg __405387_405387;
   reg _405388_405388 ; 
   reg __405388_405388;
   reg _405389_405389 ; 
   reg __405389_405389;
   reg _405390_405390 ; 
   reg __405390_405390;
   reg _405391_405391 ; 
   reg __405391_405391;
   reg _405392_405392 ; 
   reg __405392_405392;
   reg _405393_405393 ; 
   reg __405393_405393;
   reg _405394_405394 ; 
   reg __405394_405394;
   reg _405395_405395 ; 
   reg __405395_405395;
   reg _405396_405396 ; 
   reg __405396_405396;
   reg _405397_405397 ; 
   reg __405397_405397;
   reg _405398_405398 ; 
   reg __405398_405398;
   reg _405399_405399 ; 
   reg __405399_405399;
   reg _405400_405400 ; 
   reg __405400_405400;
   reg _405401_405401 ; 
   reg __405401_405401;
   reg _405402_405402 ; 
   reg __405402_405402;
   reg _405403_405403 ; 
   reg __405403_405403;
   reg _405404_405404 ; 
   reg __405404_405404;
   reg _405405_405405 ; 
   reg __405405_405405;
   reg _405406_405406 ; 
   reg __405406_405406;
   reg _405407_405407 ; 
   reg __405407_405407;
   reg _405408_405408 ; 
   reg __405408_405408;
   reg _405409_405409 ; 
   reg __405409_405409;
   reg _405410_405410 ; 
   reg __405410_405410;
   reg _405411_405411 ; 
   reg __405411_405411;
   reg _405412_405412 ; 
   reg __405412_405412;
   reg _405413_405413 ; 
   reg __405413_405413;
   reg _405414_405414 ; 
   reg __405414_405414;
   reg _405415_405415 ; 
   reg __405415_405415;
   reg _405416_405416 ; 
   reg __405416_405416;
   reg _405417_405417 ; 
   reg __405417_405417;
   reg _405418_405418 ; 
   reg __405418_405418;
   reg _405419_405419 ; 
   reg __405419_405419;
   reg _405420_405420 ; 
   reg __405420_405420;
   reg _405421_405421 ; 
   reg __405421_405421;
   reg _405422_405422 ; 
   reg __405422_405422;
   reg _405423_405423 ; 
   reg __405423_405423;
   reg _405424_405424 ; 
   reg __405424_405424;
   reg _405425_405425 ; 
   reg __405425_405425;
   reg _405426_405426 ; 
   reg __405426_405426;
   reg _405427_405427 ; 
   reg __405427_405427;
   reg _405428_405428 ; 
   reg __405428_405428;
   reg _405429_405429 ; 
   reg __405429_405429;
   reg _405430_405430 ; 
   reg __405430_405430;
   reg _405431_405431 ; 
   reg __405431_405431;
   reg _405432_405432 ; 
   reg __405432_405432;
   reg _405433_405433 ; 
   reg __405433_405433;
   reg _405434_405434 ; 
   reg __405434_405434;
   reg _405435_405435 ; 
   reg __405435_405435;
   reg _405436_405436 ; 
   reg __405436_405436;
   reg _405437_405437 ; 
   reg __405437_405437;
   reg _405438_405438 ; 
   reg __405438_405438;
   reg _405439_405439 ; 
   reg __405439_405439;
   reg _405440_405440 ; 
   reg __405440_405440;
   reg _405441_405441 ; 
   reg __405441_405441;
   reg _405442_405442 ; 
   reg __405442_405442;
   reg _405443_405443 ; 
   reg __405443_405443;
   reg _405444_405444 ; 
   reg __405444_405444;
   reg _405445_405445 ; 
   reg __405445_405445;
   reg _405446_405446 ; 
   reg __405446_405446;
   reg _405447_405447 ; 
   reg __405447_405447;
   reg _405448_405448 ; 
   reg __405448_405448;
   reg _405449_405449 ; 
   reg __405449_405449;
   reg _405450_405450 ; 
   reg __405450_405450;
   reg _405451_405451 ; 
   reg __405451_405451;
   reg _405452_405452 ; 
   reg __405452_405452;
   reg _405453_405453 ; 
   reg __405453_405453;
   reg _405454_405454 ; 
   reg __405454_405454;
   reg _405455_405455 ; 
   reg __405455_405455;
   reg _405456_405456 ; 
   reg __405456_405456;
   reg _405457_405457 ; 
   reg __405457_405457;
   reg _405458_405458 ; 
   reg __405458_405458;
   reg _405459_405459 ; 
   reg __405459_405459;
   reg _405460_405460 ; 
   reg __405460_405460;
   reg _405461_405461 ; 
   reg __405461_405461;
   reg _405462_405462 ; 
   reg __405462_405462;
   reg _405463_405463 ; 
   reg __405463_405463;
   reg _405464_405464 ; 
   reg __405464_405464;
   reg _405465_405465 ; 
   reg __405465_405465;
   reg _405466_405466 ; 
   reg __405466_405466;
   reg _405467_405467 ; 
   reg __405467_405467;
   reg _405468_405468 ; 
   reg __405468_405468;
   reg _405469_405469 ; 
   reg __405469_405469;
   reg _405470_405470 ; 
   reg __405470_405470;
   reg _405471_405471 ; 
   reg __405471_405471;
   reg _405472_405472 ; 
   reg __405472_405472;
   reg _405473_405473 ; 
   reg __405473_405473;
   reg _405474_405474 ; 
   reg __405474_405474;
   reg _405475_405475 ; 
   reg __405475_405475;
   reg _405476_405476 ; 
   reg __405476_405476;
   reg _405477_405477 ; 
   reg __405477_405477;
   reg _405478_405478 ; 
   reg __405478_405478;
   reg _405479_405479 ; 
   reg __405479_405479;
   reg _405480_405480 ; 
   reg __405480_405480;
   reg _405481_405481 ; 
   reg __405481_405481;
   reg _405482_405482 ; 
   reg __405482_405482;
   reg _405483_405483 ; 
   reg __405483_405483;
   reg _405484_405484 ; 
   reg __405484_405484;
   reg _405485_405485 ; 
   reg __405485_405485;
   reg _405486_405486 ; 
   reg __405486_405486;
   reg _405487_405487 ; 
   reg __405487_405487;
   reg _405488_405488 ; 
   reg __405488_405488;
   reg _405489_405489 ; 
   reg __405489_405489;
   reg _405490_405490 ; 
   reg __405490_405490;
   reg _405491_405491 ; 
   reg __405491_405491;
   reg _405492_405492 ; 
   reg __405492_405492;
   reg _405493_405493 ; 
   reg __405493_405493;
   reg _405494_405494 ; 
   reg __405494_405494;
   reg _405495_405495 ; 
   reg __405495_405495;
   reg _405496_405496 ; 
   reg __405496_405496;
   reg _405497_405497 ; 
   reg __405497_405497;
   reg _405498_405498 ; 
   reg __405498_405498;
   reg _405499_405499 ; 
   reg __405499_405499;
   reg _405500_405500 ; 
   reg __405500_405500;
   reg _405501_405501 ; 
   reg __405501_405501;
   reg _405502_405502 ; 
   reg __405502_405502;
   reg _405503_405503 ; 
   reg __405503_405503;
   reg _405504_405504 ; 
   reg __405504_405504;
   reg _405505_405505 ; 
   reg __405505_405505;
   reg _405506_405506 ; 
   reg __405506_405506;
   reg _405507_405507 ; 
   reg __405507_405507;
   reg _405508_405508 ; 
   reg __405508_405508;
   reg _405509_405509 ; 
   reg __405509_405509;
   reg _405510_405510 ; 
   reg __405510_405510;
   reg _405511_405511 ; 
   reg __405511_405511;
   reg _405512_405512 ; 
   reg __405512_405512;
   reg _405513_405513 ; 
   reg __405513_405513;
   reg _405514_405514 ; 
   reg __405514_405514;
   reg _405515_405515 ; 
   reg __405515_405515;
   reg _405516_405516 ; 
   reg __405516_405516;
   reg _405517_405517 ; 
   reg __405517_405517;
   reg _405518_405518 ; 
   reg __405518_405518;
   reg _405519_405519 ; 
   reg __405519_405519;
   reg _405520_405520 ; 
   reg __405520_405520;
   reg _405521_405521 ; 
   reg __405521_405521;
   reg _405522_405522 ; 
   reg __405522_405522;
   reg _405523_405523 ; 
   reg __405523_405523;
   reg _405524_405524 ; 
   reg __405524_405524;
   reg _405525_405525 ; 
   reg __405525_405525;
   reg _405526_405526 ; 
   reg __405526_405526;
   reg _405527_405527 ; 
   reg __405527_405527;
   reg _405528_405528 ; 
   reg __405528_405528;
   reg _405529_405529 ; 
   reg __405529_405529;
   reg _405530_405530 ; 
   reg __405530_405530;
   reg _405531_405531 ; 
   reg __405531_405531;
   reg _405532_405532 ; 
   reg __405532_405532;
   reg _405533_405533 ; 
   reg __405533_405533;
   reg _405534_405534 ; 
   reg __405534_405534;
   reg _405535_405535 ; 
   reg __405535_405535;
   reg _405536_405536 ; 
   reg __405536_405536;
   reg _405537_405537 ; 
   reg __405537_405537;
   reg _405538_405538 ; 
   reg __405538_405538;
   reg _405539_405539 ; 
   reg __405539_405539;
   reg _405540_405540 ; 
   reg __405540_405540;
   reg _405541_405541 ; 
   reg __405541_405541;
   reg _405542_405542 ; 
   reg __405542_405542;
   reg _405543_405543 ; 
   reg __405543_405543;
   reg _405544_405544 ; 
   reg __405544_405544;
   reg _405545_405545 ; 
   reg __405545_405545;
   reg _405546_405546 ; 
   reg __405546_405546;
   reg _405547_405547 ; 
   reg __405547_405547;
   reg _405548_405548 ; 
   reg __405548_405548;
   reg _405549_405549 ; 
   reg __405549_405549;
   reg _405550_405550 ; 
   reg __405550_405550;
   reg _405551_405551 ; 
   reg __405551_405551;
   reg _405552_405552 ; 
   reg __405552_405552;
   reg _405553_405553 ; 
   reg __405553_405553;
   reg _405554_405554 ; 
   reg __405554_405554;
   reg _405555_405555 ; 
   reg __405555_405555;
   reg _405556_405556 ; 
   reg __405556_405556;
   reg _405557_405557 ; 
   reg __405557_405557;
   reg _405558_405558 ; 
   reg __405558_405558;
   reg _405559_405559 ; 
   reg __405559_405559;
   reg _405560_405560 ; 
   reg __405560_405560;
   reg _405561_405561 ; 
   reg __405561_405561;
   reg _405562_405562 ; 
   reg __405562_405562;
   reg _405563_405563 ; 
   reg __405563_405563;
   reg _405564_405564 ; 
   reg __405564_405564;
   reg _405565_405565 ; 
   reg __405565_405565;
   reg _405566_405566 ; 
   reg __405566_405566;
   reg _405567_405567 ; 
   reg __405567_405567;
   reg _405568_405568 ; 
   reg __405568_405568;
   reg _405569_405569 ; 
   reg __405569_405569;
   reg _405570_405570 ; 
   reg __405570_405570;
   reg _405571_405571 ; 
   reg __405571_405571;
   reg _405572_405572 ; 
   reg __405572_405572;
   reg _405573_405573 ; 
   reg __405573_405573;
   reg _405574_405574 ; 
   reg __405574_405574;
   reg _405575_405575 ; 
   reg __405575_405575;
   reg _405576_405576 ; 
   reg __405576_405576;
   reg _405577_405577 ; 
   reg __405577_405577;
   reg _405578_405578 ; 
   reg __405578_405578;
   reg _405579_405579 ; 
   reg __405579_405579;
   reg _405580_405580 ; 
   reg __405580_405580;
   reg _405581_405581 ; 
   reg __405581_405581;
   reg _405582_405582 ; 
   reg __405582_405582;
   reg _405583_405583 ; 
   reg __405583_405583;
   reg _405584_405584 ; 
   reg __405584_405584;
   reg _405585_405585 ; 
   reg __405585_405585;
   reg _405586_405586 ; 
   reg __405586_405586;
   reg _405587_405587 ; 
   reg __405587_405587;
   reg _405588_405588 ; 
   reg __405588_405588;
   reg _405589_405589 ; 
   reg __405589_405589;
   reg _405590_405590 ; 
   reg __405590_405590;
   reg _405591_405591 ; 
   reg __405591_405591;
   reg _405592_405592 ; 
   reg __405592_405592;
   reg _405593_405593 ; 
   reg __405593_405593;
   reg _405594_405594 ; 
   reg __405594_405594;
   reg _405595_405595 ; 
   reg __405595_405595;
   reg _405596_405596 ; 
   reg __405596_405596;
   reg _405597_405597 ; 
   reg __405597_405597;
   reg _405598_405598 ; 
   reg __405598_405598;
   reg _405599_405599 ; 
   reg __405599_405599;
   reg _405600_405600 ; 
   reg __405600_405600;
   reg _405601_405601 ; 
   reg __405601_405601;
   reg _405602_405602 ; 
   reg __405602_405602;
   reg _405603_405603 ; 
   reg __405603_405603;
   reg _405604_405604 ; 
   reg __405604_405604;
   reg _405605_405605 ; 
   reg __405605_405605;
   reg _405606_405606 ; 
   reg __405606_405606;
   reg _405607_405607 ; 
   reg __405607_405607;
   reg _405608_405608 ; 
   reg __405608_405608;
   reg _405609_405609 ; 
   reg __405609_405609;
   reg _405610_405610 ; 
   reg __405610_405610;
   reg _405611_405611 ; 
   reg __405611_405611;
   reg _405612_405612 ; 
   reg __405612_405612;
   reg _405613_405613 ; 
   reg __405613_405613;
   reg _405614_405614 ; 
   reg __405614_405614;
   reg _405615_405615 ; 
   reg __405615_405615;
   reg _405616_405616 ; 
   reg __405616_405616;
   reg _405617_405617 ; 
   reg __405617_405617;
   reg _405618_405618 ; 
   reg __405618_405618;
   reg _405619_405619 ; 
   reg __405619_405619;
   reg _405620_405620 ; 
   reg __405620_405620;
   reg _405621_405621 ; 
   reg __405621_405621;
   reg _405622_405622 ; 
   reg __405622_405622;
   reg _405623_405623 ; 
   reg __405623_405623;
   reg _405624_405624 ; 
   reg __405624_405624;
   reg _405625_405625 ; 
   reg __405625_405625;
   reg _405626_405626 ; 
   reg __405626_405626;
   reg _405627_405627 ; 
   reg __405627_405627;
   reg _405628_405628 ; 
   reg __405628_405628;
   reg _405629_405629 ; 
   reg __405629_405629;
   reg _405630_405630 ; 
   reg __405630_405630;
   reg _405631_405631 ; 
   reg __405631_405631;
   reg _405632_405632 ; 
   reg __405632_405632;
   reg _405633_405633 ; 
   reg __405633_405633;
   reg _405634_405634 ; 
   reg __405634_405634;
   reg _405635_405635 ; 
   reg __405635_405635;
   reg _405636_405636 ; 
   reg __405636_405636;
   reg _405637_405637 ; 
   reg __405637_405637;
   reg _405638_405638 ; 
   reg __405638_405638;
   reg _405639_405639 ; 
   reg __405639_405639;
   reg _405640_405640 ; 
   reg __405640_405640;
   reg _405641_405641 ; 
   reg __405641_405641;
   reg _405642_405642 ; 
   reg __405642_405642;
   reg _405643_405643 ; 
   reg __405643_405643;
   reg _405644_405644 ; 
   reg __405644_405644;
   reg _405645_405645 ; 
   reg __405645_405645;
   reg _405646_405646 ; 
   reg __405646_405646;
   reg _405647_405647 ; 
   reg __405647_405647;
   reg _405648_405648 ; 
   reg __405648_405648;
   reg _405649_405649 ; 
   reg __405649_405649;
   reg _405650_405650 ; 
   reg __405650_405650;
   reg _405651_405651 ; 
   reg __405651_405651;
   reg _405652_405652 ; 
   reg __405652_405652;
   reg _405653_405653 ; 
   reg __405653_405653;
   reg _405654_405654 ; 
   reg __405654_405654;
   reg _405655_405655 ; 
   reg __405655_405655;
   reg _405656_405656 ; 
   reg __405656_405656;
   reg _405657_405657 ; 
   reg __405657_405657;
   reg _405658_405658 ; 
   reg __405658_405658;
   reg _405659_405659 ; 
   reg __405659_405659;
   reg _405660_405660 ; 
   reg __405660_405660;
   reg _405661_405661 ; 
   reg __405661_405661;
   reg _405662_405662 ; 
   reg __405662_405662;
   reg _405663_405663 ; 
   reg __405663_405663;
   reg _405664_405664 ; 
   reg __405664_405664;
   reg _405665_405665 ; 
   reg __405665_405665;
   reg _405666_405666 ; 
   reg __405666_405666;
   reg _405667_405667 ; 
   reg __405667_405667;
   reg _405668_405668 ; 
   reg __405668_405668;
   reg _405669_405669 ; 
   reg __405669_405669;
   reg _405670_405670 ; 
   reg __405670_405670;
   reg _405671_405671 ; 
   reg __405671_405671;
   reg _405672_405672 ; 
   reg __405672_405672;
   reg _405673_405673 ; 
   reg __405673_405673;
   reg _405674_405674 ; 
   reg __405674_405674;
   reg _405675_405675 ; 
   reg __405675_405675;
   reg _405676_405676 ; 
   reg __405676_405676;
   reg _405677_405677 ; 
   reg __405677_405677;
   reg _405678_405678 ; 
   reg __405678_405678;
   reg _405679_405679 ; 
   reg __405679_405679;
   reg _405680_405680 ; 
   reg __405680_405680;
   reg _405681_405681 ; 
   reg __405681_405681;
   reg _405682_405682 ; 
   reg __405682_405682;
   reg _405683_405683 ; 
   reg __405683_405683;
   reg _405684_405684 ; 
   reg __405684_405684;
   reg _405685_405685 ; 
   reg __405685_405685;
   reg _405686_405686 ; 
   reg __405686_405686;
   reg _405687_405687 ; 
   reg __405687_405687;
   reg _405688_405688 ; 
   reg __405688_405688;
   reg _405689_405689 ; 
   reg __405689_405689;
   reg _405690_405690 ; 
   reg __405690_405690;
   reg _405691_405691 ; 
   reg __405691_405691;
   reg _405692_405692 ; 
   reg __405692_405692;
   reg _405693_405693 ; 
   reg __405693_405693;
   reg _405694_405694 ; 
   reg __405694_405694;
   reg _405695_405695 ; 
   reg __405695_405695;
   reg _405696_405696 ; 
   reg __405696_405696;
   reg _405697_405697 ; 
   reg __405697_405697;
   reg _405698_405698 ; 
   reg __405698_405698;
   reg _405699_405699 ; 
   reg __405699_405699;
   reg _405700_405700 ; 
   reg __405700_405700;
   reg _405701_405701 ; 
   reg __405701_405701;
   reg _405702_405702 ; 
   reg __405702_405702;
   reg _405703_405703 ; 
   reg __405703_405703;
   reg _405704_405704 ; 
   reg __405704_405704;
   reg _405705_405705 ; 
   reg __405705_405705;
   reg _405706_405706 ; 
   reg __405706_405706;
   reg _405707_405707 ; 
   reg __405707_405707;
   reg _405708_405708 ; 
   reg __405708_405708;
   reg _405709_405709 ; 
   reg __405709_405709;
   reg _405710_405710 ; 
   reg __405710_405710;
   reg _405711_405711 ; 
   reg __405711_405711;
   reg _405712_405712 ; 
   reg __405712_405712;
   reg _405713_405713 ; 
   reg __405713_405713;
   reg _405714_405714 ; 
   reg __405714_405714;
   reg _405715_405715 ; 
   reg __405715_405715;
   reg _405716_405716 ; 
   reg __405716_405716;
   reg _405717_405717 ; 
   reg __405717_405717;
   reg _405718_405718 ; 
   reg __405718_405718;
   reg _405719_405719 ; 
   reg __405719_405719;
   reg _405720_405720 ; 
   reg __405720_405720;
   reg _405721_405721 ; 
   reg __405721_405721;
   reg _405722_405722 ; 
   reg __405722_405722;
   reg _405723_405723 ; 
   reg __405723_405723;
   reg _405724_405724 ; 
   reg __405724_405724;
   reg _405725_405725 ; 
   reg __405725_405725;
   reg _405726_405726 ; 
   reg __405726_405726;
   reg _405727_405727 ; 
   reg __405727_405727;
   reg _405728_405728 ; 
   reg __405728_405728;
   reg _405729_405729 ; 
   reg __405729_405729;
   reg _405730_405730 ; 
   reg __405730_405730;
   reg _405731_405731 ; 
   reg __405731_405731;
   reg _405732_405732 ; 
   reg __405732_405732;
   reg _405733_405733 ; 
   reg __405733_405733;
   reg _405734_405734 ; 
   reg __405734_405734;
   reg _405735_405735 ; 
   reg __405735_405735;
   reg _405736_405736 ; 
   reg __405736_405736;
   reg _405737_405737 ; 
   reg __405737_405737;
   reg _405738_405738 ; 
   reg __405738_405738;
   reg _405739_405739 ; 
   reg __405739_405739;
   reg _405740_405740 ; 
   reg __405740_405740;
   reg _405741_405741 ; 
   reg __405741_405741;
   reg _405742_405742 ; 
   reg __405742_405742;
   reg _405743_405743 ; 
   reg __405743_405743;
   reg _405744_405744 ; 
   reg __405744_405744;
   reg _405745_405745 ; 
   reg __405745_405745;
   reg _405746_405746 ; 
   reg __405746_405746;
   reg _405747_405747 ; 
   reg __405747_405747;
   reg _405748_405748 ; 
   reg __405748_405748;
   reg _405749_405749 ; 
   reg __405749_405749;
   reg _405750_405750 ; 
   reg __405750_405750;
   reg _405751_405751 ; 
   reg __405751_405751;
   reg _405752_405752 ; 
   reg __405752_405752;
   reg _405753_405753 ; 
   reg __405753_405753;
   reg _405754_405754 ; 
   reg __405754_405754;
   reg _405755_405755 ; 
   reg __405755_405755;
   reg _405756_405756 ; 
   reg __405756_405756;
   reg _405757_405757 ; 
   reg __405757_405757;
   reg _405758_405758 ; 
   reg __405758_405758;
   reg _405759_405759 ; 
   reg __405759_405759;
   reg _405760_405760 ; 
   reg __405760_405760;
   reg _405761_405761 ; 
   reg __405761_405761;
   reg _405762_405762 ; 
   reg __405762_405762;
   reg _405763_405763 ; 
   reg __405763_405763;
   reg _405764_405764 ; 
   reg __405764_405764;
   reg _405765_405765 ; 
   reg __405765_405765;
   reg _405766_405766 ; 
   reg __405766_405766;
   reg _405767_405767 ; 
   reg __405767_405767;
   reg _405768_405768 ; 
   reg __405768_405768;
   reg _405769_405769 ; 
   reg __405769_405769;
   reg _405770_405770 ; 
   reg __405770_405770;
   reg _405771_405771 ; 
   reg __405771_405771;
   reg _405772_405772 ; 
   reg __405772_405772;
   reg _405773_405773 ; 
   reg __405773_405773;
   reg _405774_405774 ; 
   reg __405774_405774;
   reg _405775_405775 ; 
   reg __405775_405775;
   reg _405776_405776 ; 
   reg __405776_405776;
   reg _405777_405777 ; 
   reg __405777_405777;
   reg _405778_405778 ; 
   reg __405778_405778;
   reg _405779_405779 ; 
   reg __405779_405779;
   reg _405780_405780 ; 
   reg __405780_405780;
   reg _405781_405781 ; 
   reg __405781_405781;
   reg _405782_405782 ; 
   reg __405782_405782;
   reg _405783_405783 ; 
   reg __405783_405783;
   reg _405784_405784 ; 
   reg __405784_405784;
   reg _405785_405785 ; 
   reg __405785_405785;
   reg _405786_405786 ; 
   reg __405786_405786;
   reg _405787_405787 ; 
   reg __405787_405787;
   reg _405788_405788 ; 
   reg __405788_405788;
   reg _405789_405789 ; 
   reg __405789_405789;
   reg _405790_405790 ; 
   reg __405790_405790;
   reg _405791_405791 ; 
   reg __405791_405791;
   reg _405792_405792 ; 
   reg __405792_405792;
   reg _405793_405793 ; 
   reg __405793_405793;
   reg _405794_405794 ; 
   reg __405794_405794;
   reg _405795_405795 ; 
   reg __405795_405795;
   reg _405796_405796 ; 
   reg __405796_405796;
   reg _405797_405797 ; 
   reg __405797_405797;
   reg _405798_405798 ; 
   reg __405798_405798;
   reg _405799_405799 ; 
   reg __405799_405799;
   reg _405800_405800 ; 
   reg __405800_405800;
   reg _405801_405801 ; 
   reg __405801_405801;
   reg _405802_405802 ; 
   reg __405802_405802;
   reg _405803_405803 ; 
   reg __405803_405803;
   reg _405804_405804 ; 
   reg __405804_405804;
   reg _405805_405805 ; 
   reg __405805_405805;
   reg _405806_405806 ; 
   reg __405806_405806;
   reg _405807_405807 ; 
   reg __405807_405807;
   reg _405808_405808 ; 
   reg __405808_405808;
   reg _405809_405809 ; 
   reg __405809_405809;
   reg _405810_405810 ; 
   reg __405810_405810;
   reg _405811_405811 ; 
   reg __405811_405811;
   reg _405812_405812 ; 
   reg __405812_405812;
   reg _405813_405813 ; 
   reg __405813_405813;
   reg _405814_405814 ; 
   reg __405814_405814;
   reg _405815_405815 ; 
   reg __405815_405815;
   reg _405816_405816 ; 
   reg __405816_405816;
   reg _405817_405817 ; 
   reg __405817_405817;
   reg _405818_405818 ; 
   reg __405818_405818;
   reg _405819_405819 ; 
   reg __405819_405819;
   reg _405820_405820 ; 
   reg __405820_405820;
   reg _405821_405821 ; 
   reg __405821_405821;
   reg _405822_405822 ; 
   reg __405822_405822;
   reg _405823_405823 ; 
   reg __405823_405823;
   reg _405824_405824 ; 
   reg __405824_405824;
   reg _405825_405825 ; 
   reg __405825_405825;
   reg _405826_405826 ; 
   reg __405826_405826;
   reg _405827_405827 ; 
   reg __405827_405827;
   reg _405828_405828 ; 
   reg __405828_405828;
   reg _405829_405829 ; 
   reg __405829_405829;
   reg _405830_405830 ; 
   reg __405830_405830;
   reg _405831_405831 ; 
   reg __405831_405831;
   reg _405832_405832 ; 
   reg __405832_405832;
   reg _405833_405833 ; 
   reg __405833_405833;
   reg _405834_405834 ; 
   reg __405834_405834;
   reg _405835_405835 ; 
   reg __405835_405835;
   reg _405836_405836 ; 
   reg __405836_405836;
   reg _405837_405837 ; 
   reg __405837_405837;
   reg _405838_405838 ; 
   reg __405838_405838;
   reg _405839_405839 ; 
   reg __405839_405839;
   reg _405840_405840 ; 
   reg __405840_405840;
   reg _405841_405841 ; 
   reg __405841_405841;
   reg _405842_405842 ; 
   reg __405842_405842;
   reg _405843_405843 ; 
   reg __405843_405843;
   reg _405844_405844 ; 
   reg __405844_405844;
   reg _405845_405845 ; 
   reg __405845_405845;
   reg _405846_405846 ; 
   reg __405846_405846;
   reg _405847_405847 ; 
   reg __405847_405847;
   reg _405848_405848 ; 
   reg __405848_405848;
   reg _405849_405849 ; 
   reg __405849_405849;
   reg _405850_405850 ; 
   reg __405850_405850;
   reg _405851_405851 ; 
   reg __405851_405851;
   reg _405852_405852 ; 
   reg __405852_405852;
   reg _405853_405853 ; 
   reg __405853_405853;
   reg _405854_405854 ; 
   reg __405854_405854;
   reg _405855_405855 ; 
   reg __405855_405855;
   reg _405856_405856 ; 
   reg __405856_405856;
   reg _405857_405857 ; 
   reg __405857_405857;
   reg _405858_405858 ; 
   reg __405858_405858;
   reg _405859_405859 ; 
   reg __405859_405859;
   reg _405860_405860 ; 
   reg __405860_405860;
   reg _405861_405861 ; 
   reg __405861_405861;
   reg _405862_405862 ; 
   reg __405862_405862;
   reg _405863_405863 ; 
   reg __405863_405863;
   reg _405864_405864 ; 
   reg __405864_405864;
   reg _405865_405865 ; 
   reg __405865_405865;
   reg _405866_405866 ; 
   reg __405866_405866;
   reg _405867_405867 ; 
   reg __405867_405867;
   reg _405868_405868 ; 
   reg __405868_405868;
   reg _405869_405869 ; 
   reg __405869_405869;
   reg _405870_405870 ; 
   reg __405870_405870;
   reg _405871_405871 ; 
   reg __405871_405871;
   reg _405872_405872 ; 
   reg __405872_405872;
   reg _405873_405873 ; 
   reg __405873_405873;
   reg _405874_405874 ; 
   reg __405874_405874;
   reg _405875_405875 ; 
   reg __405875_405875;
   reg _405876_405876 ; 
   reg __405876_405876;
   reg _405877_405877 ; 
   reg __405877_405877;
   reg _405878_405878 ; 
   reg __405878_405878;
   reg _405879_405879 ; 
   reg __405879_405879;
   reg _405880_405880 ; 
   reg __405880_405880;
   reg _405881_405881 ; 
   reg __405881_405881;
   reg _405882_405882 ; 
   reg __405882_405882;
   reg _405883_405883 ; 
   reg __405883_405883;
   reg _405884_405884 ; 
   reg __405884_405884;
   reg _405885_405885 ; 
   reg __405885_405885;
   reg _405886_405886 ; 
   reg __405886_405886;
   reg _405887_405887 ; 
   reg __405887_405887;
   reg _405888_405888 ; 
   reg __405888_405888;
   reg _405889_405889 ; 
   reg __405889_405889;
   reg _405890_405890 ; 
   reg __405890_405890;
   reg _405891_405891 ; 
   reg __405891_405891;
   reg _405892_405892 ; 
   reg __405892_405892;
   reg _405893_405893 ; 
   reg __405893_405893;
   reg _405894_405894 ; 
   reg __405894_405894;
   reg _405895_405895 ; 
   reg __405895_405895;
   reg _405896_405896 ; 
   reg __405896_405896;
   reg _405897_405897 ; 
   reg __405897_405897;
   reg _405898_405898 ; 
   reg __405898_405898;
   reg _405899_405899 ; 
   reg __405899_405899;
   reg _405900_405900 ; 
   reg __405900_405900;
   reg _405901_405901 ; 
   reg __405901_405901;
   reg _405902_405902 ; 
   reg __405902_405902;
   reg _405903_405903 ; 
   reg __405903_405903;
   reg _405904_405904 ; 
   reg __405904_405904;
   reg _405905_405905 ; 
   reg __405905_405905;
   reg _405906_405906 ; 
   reg __405906_405906;
   reg _405907_405907 ; 
   reg __405907_405907;
   reg _405908_405908 ; 
   reg __405908_405908;
   reg _405909_405909 ; 
   reg __405909_405909;
   reg _405910_405910 ; 
   reg __405910_405910;
   reg _405911_405911 ; 
   reg __405911_405911;
   reg _405912_405912 ; 
   reg __405912_405912;
   reg _405913_405913 ; 
   reg __405913_405913;
   reg _405914_405914 ; 
   reg __405914_405914;
   reg _405915_405915 ; 
   reg __405915_405915;
   reg _405916_405916 ; 
   reg __405916_405916;
   reg _405917_405917 ; 
   reg __405917_405917;
   reg _405918_405918 ; 
   reg __405918_405918;
   reg _405919_405919 ; 
   reg __405919_405919;
   reg _405920_405920 ; 
   reg __405920_405920;
   reg _405921_405921 ; 
   reg __405921_405921;
   reg _405922_405922 ; 
   reg __405922_405922;
   reg _405923_405923 ; 
   reg __405923_405923;
   reg _405924_405924 ; 
   reg __405924_405924;
   reg _405925_405925 ; 
   reg __405925_405925;
   reg _405926_405926 ; 
   reg __405926_405926;
   reg _405927_405927 ; 
   reg __405927_405927;
   reg _405928_405928 ; 
   reg __405928_405928;
   reg _405929_405929 ; 
   reg __405929_405929;
   reg _405930_405930 ; 
   reg __405930_405930;
   reg _405931_405931 ; 
   reg __405931_405931;
   reg _405932_405932 ; 
   reg __405932_405932;
   reg _405933_405933 ; 
   reg __405933_405933;
   reg _405934_405934 ; 
   reg __405934_405934;
   reg _405935_405935 ; 
   reg __405935_405935;
   reg _405936_405936 ; 
   reg __405936_405936;
   reg _405937_405937 ; 
   reg __405937_405937;
   reg _405938_405938 ; 
   reg __405938_405938;
   reg _405939_405939 ; 
   reg __405939_405939;
   reg _405940_405940 ; 
   reg __405940_405940;
   reg _405941_405941 ; 
   reg __405941_405941;
   reg _405942_405942 ; 
   reg __405942_405942;
   reg _405943_405943 ; 
   reg __405943_405943;
   reg _405944_405944 ; 
   reg __405944_405944;
   reg _405945_405945 ; 
   reg __405945_405945;
   reg _405946_405946 ; 
   reg __405946_405946;
   reg _405947_405947 ; 
   reg __405947_405947;
   reg _405948_405948 ; 
   reg __405948_405948;
   reg _405949_405949 ; 
   reg __405949_405949;
   reg _405950_405950 ; 
   reg __405950_405950;
   reg _405951_405951 ; 
   reg __405951_405951;
   reg _405952_405952 ; 
   reg __405952_405952;
   reg _405953_405953 ; 
   reg __405953_405953;
   reg _405954_405954 ; 
   reg __405954_405954;
   reg _405955_405955 ; 
   reg __405955_405955;
   reg _405956_405956 ; 
   reg __405956_405956;
   reg _405957_405957 ; 
   reg __405957_405957;
   reg _405958_405958 ; 
   reg __405958_405958;
   reg _405959_405959 ; 
   reg __405959_405959;
   reg _405960_405960 ; 
   reg __405960_405960;
   reg _405961_405961 ; 
   reg __405961_405961;
   reg _405962_405962 ; 
   reg __405962_405962;
   reg _405963_405963 ; 
   reg __405963_405963;
   reg _405964_405964 ; 
   reg __405964_405964;
   reg _405965_405965 ; 
   reg __405965_405965;
   reg _405966_405966 ; 
   reg __405966_405966;
   reg _405967_405967 ; 
   reg __405967_405967;
   reg _405968_405968 ; 
   reg __405968_405968;
   reg _405969_405969 ; 
   reg __405969_405969;
   reg _405970_405970 ; 
   reg __405970_405970;
   reg _405971_405971 ; 
   reg __405971_405971;
   reg _405972_405972 ; 
   reg __405972_405972;
   reg _405973_405973 ; 
   reg __405973_405973;
   reg _405974_405974 ; 
   reg __405974_405974;
   reg _405975_405975 ; 
   reg __405975_405975;
   reg _405976_405976 ; 
   reg __405976_405976;
   reg _405977_405977 ; 
   reg __405977_405977;
   reg _405978_405978 ; 
   reg __405978_405978;
   reg _405979_405979 ; 
   reg __405979_405979;
   reg _405980_405980 ; 
   reg __405980_405980;
   reg _405981_405981 ; 
   reg __405981_405981;
   reg _405982_405982 ; 
   reg __405982_405982;
   reg _405983_405983 ; 
   reg __405983_405983;
   reg _405984_405984 ; 
   reg __405984_405984;
   reg _405985_405985 ; 
   reg __405985_405985;
   reg _405986_405986 ; 
   reg __405986_405986;
   reg _405987_405987 ; 
   reg __405987_405987;
   reg _405988_405988 ; 
   reg __405988_405988;
   reg _405989_405989 ; 
   reg __405989_405989;
   reg _405990_405990 ; 
   reg __405990_405990;
   reg _405991_405991 ; 
   reg __405991_405991;
   reg _405992_405992 ; 
   reg __405992_405992;
   reg _405993_405993 ; 
   reg __405993_405993;
   reg _405994_405994 ; 
   reg __405994_405994;
   reg _405995_405995 ; 
   reg __405995_405995;
   reg _405996_405996 ; 
   reg __405996_405996;
   reg _405997_405997 ; 
   reg __405997_405997;
   reg _405998_405998 ; 
   reg __405998_405998;
   reg _405999_405999 ; 
   reg __405999_405999;
   reg _406000_406000 ; 
   reg __406000_406000;
   reg _406001_406001 ; 
   reg __406001_406001;
   reg _406002_406002 ; 
   reg __406002_406002;
   reg _406003_406003 ; 
   reg __406003_406003;
   reg _406004_406004 ; 
   reg __406004_406004;
   reg _406005_406005 ; 
   reg __406005_406005;
   reg _406006_406006 ; 
   reg __406006_406006;
   reg _406007_406007 ; 
   reg __406007_406007;
   reg _406008_406008 ; 
   reg __406008_406008;
   reg _406009_406009 ; 
   reg __406009_406009;
   reg _406010_406010 ; 
   reg __406010_406010;
   reg _406011_406011 ; 
   reg __406011_406011;
   reg _406012_406012 ; 
   reg __406012_406012;
   reg _406013_406013 ; 
   reg __406013_406013;
   reg _406014_406014 ; 
   reg __406014_406014;
   reg _406015_406015 ; 
   reg __406015_406015;
   reg _406016_406016 ; 
   reg __406016_406016;
   reg _406017_406017 ; 
   reg __406017_406017;
   reg _406018_406018 ; 
   reg __406018_406018;
   reg _406019_406019 ; 
   reg __406019_406019;
   reg _406020_406020 ; 
   reg __406020_406020;
   reg _406021_406021 ; 
   reg __406021_406021;
   reg _406022_406022 ; 
   reg __406022_406022;
   reg _406023_406023 ; 
   reg __406023_406023;
   reg _406024_406024 ; 
   reg __406024_406024;
   reg _406025_406025 ; 
   reg __406025_406025;
   reg _406026_406026 ; 
   reg __406026_406026;
   reg _406027_406027 ; 
   reg __406027_406027;
   reg _406028_406028 ; 
   reg __406028_406028;
   reg _406029_406029 ; 
   reg __406029_406029;
   reg _406030_406030 ; 
   reg __406030_406030;
   reg _406031_406031 ; 
   reg __406031_406031;
   reg _406032_406032 ; 
   reg __406032_406032;
   reg _406033_406033 ; 
   reg __406033_406033;
   reg _406034_406034 ; 
   reg __406034_406034;
   reg _406035_406035 ; 
   reg __406035_406035;
   reg _406036_406036 ; 
   reg __406036_406036;
   reg _406037_406037 ; 
   reg __406037_406037;
   reg _406038_406038 ; 
   reg __406038_406038;
   reg _406039_406039 ; 
   reg __406039_406039;
   reg _406040_406040 ; 
   reg __406040_406040;
   reg _406041_406041 ; 
   reg __406041_406041;
   reg _406042_406042 ; 
   reg __406042_406042;
   reg _406043_406043 ; 
   reg __406043_406043;
   reg _406044_406044 ; 
   reg __406044_406044;
   reg _406045_406045 ; 
   reg __406045_406045;
   reg _406046_406046 ; 
   reg __406046_406046;
   reg _406047_406047 ; 
   reg __406047_406047;
   reg _406048_406048 ; 
   reg __406048_406048;
   reg _406049_406049 ; 
   reg __406049_406049;
   reg _406050_406050 ; 
   reg __406050_406050;
   reg _406051_406051 ; 
   reg __406051_406051;
   reg _406052_406052 ; 
   reg __406052_406052;
   reg _406053_406053 ; 
   reg __406053_406053;
   reg _406054_406054 ; 
   reg __406054_406054;
   reg _406055_406055 ; 
   reg __406055_406055;
   reg _406056_406056 ; 
   reg __406056_406056;
   reg _406057_406057 ; 
   reg __406057_406057;
   reg _406058_406058 ; 
   reg __406058_406058;
   reg _406059_406059 ; 
   reg __406059_406059;
   reg _406060_406060 ; 
   reg __406060_406060;
   reg _406061_406061 ; 
   reg __406061_406061;
   reg _406062_406062 ; 
   reg __406062_406062;
   reg _406063_406063 ; 
   reg __406063_406063;
   reg _406064_406064 ; 
   reg __406064_406064;
   reg _406065_406065 ; 
   reg __406065_406065;
   reg _406066_406066 ; 
   reg __406066_406066;
   reg _406067_406067 ; 
   reg __406067_406067;
   reg _406068_406068 ; 
   reg __406068_406068;
   reg _406069_406069 ; 
   reg __406069_406069;
   reg _406070_406070 ; 
   reg __406070_406070;
   reg _406071_406071 ; 
   reg __406071_406071;
   reg _406072_406072 ; 
   reg __406072_406072;
   reg _406073_406073 ; 
   reg __406073_406073;
   reg _406074_406074 ; 
   reg __406074_406074;
   reg _406075_406075 ; 
   reg __406075_406075;
   reg _406076_406076 ; 
   reg __406076_406076;
   reg _406077_406077 ; 
   reg __406077_406077;
   reg _406078_406078 ; 
   reg __406078_406078;
   reg _406079_406079 ; 
   reg __406079_406079;
   reg _406080_406080 ; 
   reg __406080_406080;
   reg _406081_406081 ; 
   reg __406081_406081;
   reg _406082_406082 ; 
   reg __406082_406082;
   reg _406083_406083 ; 
   reg __406083_406083;
   reg _406084_406084 ; 
   reg __406084_406084;
   reg _406085_406085 ; 
   reg __406085_406085;
   reg _406086_406086 ; 
   reg __406086_406086;
   reg _406087_406087 ; 
   reg __406087_406087;
   reg _406088_406088 ; 
   reg __406088_406088;
   reg _406089_406089 ; 
   reg __406089_406089;
   reg _406090_406090 ; 
   reg __406090_406090;
   reg _406091_406091 ; 
   reg __406091_406091;
   reg _406092_406092 ; 
   reg __406092_406092;
   reg _406093_406093 ; 
   reg __406093_406093;
   reg _406094_406094 ; 
   reg __406094_406094;
   reg _406095_406095 ; 
   reg __406095_406095;
   reg _406096_406096 ; 
   reg __406096_406096;
   reg _406097_406097 ; 
   reg __406097_406097;
   reg _406098_406098 ; 
   reg __406098_406098;
   reg _406099_406099 ; 
   reg __406099_406099;
   reg _406100_406100 ; 
   reg __406100_406100;
   reg _406101_406101 ; 
   reg __406101_406101;
   reg _406102_406102 ; 
   reg __406102_406102;
   reg _406103_406103 ; 
   reg __406103_406103;
   reg _406104_406104 ; 
   reg __406104_406104;
   reg _406105_406105 ; 
   reg __406105_406105;
   reg _406106_406106 ; 
   reg __406106_406106;
   reg _406107_406107 ; 
   reg __406107_406107;
   reg _406108_406108 ; 
   reg __406108_406108;
   reg _406109_406109 ; 
   reg __406109_406109;
   reg _406110_406110 ; 
   reg __406110_406110;
   reg _406111_406111 ; 
   reg __406111_406111;
   reg _406112_406112 ; 
   reg __406112_406112;
   reg _406113_406113 ; 
   reg __406113_406113;
   reg _406114_406114 ; 
   reg __406114_406114;
   reg _406115_406115 ; 
   reg __406115_406115;
   reg _406116_406116 ; 
   reg __406116_406116;
   reg _406117_406117 ; 
   reg __406117_406117;
   reg _406118_406118 ; 
   reg __406118_406118;
   reg _406119_406119 ; 
   reg __406119_406119;
   reg _406120_406120 ; 
   reg __406120_406120;
   reg _406121_406121 ; 
   reg __406121_406121;
   reg _406122_406122 ; 
   reg __406122_406122;
   reg _406123_406123 ; 
   reg __406123_406123;
   reg _406124_406124 ; 
   reg __406124_406124;
   reg _406125_406125 ; 
   reg __406125_406125;
   reg _406126_406126 ; 
   reg __406126_406126;
   reg _406127_406127 ; 
   reg __406127_406127;
   reg _406128_406128 ; 
   reg __406128_406128;
   reg _406129_406129 ; 
   reg __406129_406129;
   reg _406130_406130 ; 
   reg __406130_406130;
   reg _406131_406131 ; 
   reg __406131_406131;
   reg _406132_406132 ; 
   reg __406132_406132;
   reg _406133_406133 ; 
   reg __406133_406133;
   reg _406134_406134 ; 
   reg __406134_406134;
   reg _406135_406135 ; 
   reg __406135_406135;
   reg _406136_406136 ; 
   reg __406136_406136;
   reg _406137_406137 ; 
   reg __406137_406137;
   reg _406138_406138 ; 
   reg __406138_406138;
   reg _406139_406139 ; 
   reg __406139_406139;
   reg _406140_406140 ; 
   reg __406140_406140;
   reg _406141_406141 ; 
   reg __406141_406141;
   reg _406142_406142 ; 
   reg __406142_406142;
   reg _406143_406143 ; 
   reg __406143_406143;
   reg _406144_406144 ; 
   reg __406144_406144;
   reg _406145_406145 ; 
   reg __406145_406145;
   reg _406146_406146 ; 
   reg __406146_406146;
   reg _406147_406147 ; 
   reg __406147_406147;
   reg _406148_406148 ; 
   reg __406148_406148;
   reg _406149_406149 ; 
   reg __406149_406149;
   reg _406150_406150 ; 
   reg __406150_406150;
   reg _406151_406151 ; 
   reg __406151_406151;
   reg _406152_406152 ; 
   reg __406152_406152;
   reg _406153_406153 ; 
   reg __406153_406153;
   reg _406154_406154 ; 
   reg __406154_406154;
   reg _406155_406155 ; 
   reg __406155_406155;
   reg _406156_406156 ; 
   reg __406156_406156;
   reg _406157_406157 ; 
   reg __406157_406157;
   reg _406158_406158 ; 
   reg __406158_406158;
   reg _406159_406159 ; 
   reg __406159_406159;
   reg _406160_406160 ; 
   reg __406160_406160;
   reg _406161_406161 ; 
   reg __406161_406161;
   reg _406162_406162 ; 
   reg __406162_406162;
   reg _406163_406163 ; 
   reg __406163_406163;
   reg _406164_406164 ; 
   reg __406164_406164;
   reg _406165_406165 ; 
   reg __406165_406165;
   reg _406166_406166 ; 
   reg __406166_406166;
   reg _406167_406167 ; 
   reg __406167_406167;
   reg _406168_406168 ; 
   reg __406168_406168;
   reg _406169_406169 ; 
   reg __406169_406169;
   reg _406170_406170 ; 
   reg __406170_406170;
   reg _406171_406171 ; 
   reg __406171_406171;
   reg _406172_406172 ; 
   reg __406172_406172;
   reg _406173_406173 ; 
   reg __406173_406173;
   reg _406174_406174 ; 
   reg __406174_406174;
   reg _406175_406175 ; 
   reg __406175_406175;
   reg _406176_406176 ; 
   reg __406176_406176;
   reg _406177_406177 ; 
   reg __406177_406177;
   reg _406178_406178 ; 
   reg __406178_406178;
   reg _406179_406179 ; 
   reg __406179_406179;
   reg _406180_406180 ; 
   reg __406180_406180;
   reg _406181_406181 ; 
   reg __406181_406181;
   reg _406182_406182 ; 
   reg __406182_406182;
   reg _406183_406183 ; 
   reg __406183_406183;
   reg _406184_406184 ; 
   reg __406184_406184;
   reg _406185_406185 ; 
   reg __406185_406185;
   reg _406186_406186 ; 
   reg __406186_406186;
   reg _406187_406187 ; 
   reg __406187_406187;
   reg _406188_406188 ; 
   reg __406188_406188;
   reg _406189_406189 ; 
   reg __406189_406189;
   reg _406190_406190 ; 
   reg __406190_406190;
   reg _406191_406191 ; 
   reg __406191_406191;
   reg _406192_406192 ; 
   reg __406192_406192;
   reg _406193_406193 ; 
   reg __406193_406193;
   reg _406194_406194 ; 
   reg __406194_406194;
   reg _406195_406195 ; 
   reg __406195_406195;
   reg _406196_406196 ; 
   reg __406196_406196;
   reg _406197_406197 ; 
   reg __406197_406197;
   reg _406198_406198 ; 
   reg __406198_406198;
   reg _406199_406199 ; 
   reg __406199_406199;
   reg _406200_406200 ; 
   reg __406200_406200;
   reg _406201_406201 ; 
   reg __406201_406201;
   reg _406202_406202 ; 
   reg __406202_406202;
   reg _406203_406203 ; 
   reg __406203_406203;
   reg _406204_406204 ; 
   reg __406204_406204;
   reg _406205_406205 ; 
   reg __406205_406205;
   reg _406206_406206 ; 
   reg __406206_406206;
   reg _406207_406207 ; 
   reg __406207_406207;
   reg _406208_406208 ; 
   reg __406208_406208;
   reg _406209_406209 ; 
   reg __406209_406209;
   reg _406210_406210 ; 
   reg __406210_406210;
   reg _406211_406211 ; 
   reg __406211_406211;
   reg _406212_406212 ; 
   reg __406212_406212;
   reg _406213_406213 ; 
   reg __406213_406213;
   reg _406214_406214 ; 
   reg __406214_406214;
   reg _406215_406215 ; 
   reg __406215_406215;
   reg _406216_406216 ; 
   reg __406216_406216;
   reg _406217_406217 ; 
   reg __406217_406217;
   reg _406218_406218 ; 
   reg __406218_406218;
   reg _406219_406219 ; 
   reg __406219_406219;
   reg _406220_406220 ; 
   reg __406220_406220;
   reg _406221_406221 ; 
   reg __406221_406221;
   reg _406222_406222 ; 
   reg __406222_406222;
   reg _406223_406223 ; 
   reg __406223_406223;
   reg _406224_406224 ; 
   reg __406224_406224;
   reg _406225_406225 ; 
   reg __406225_406225;
   reg _406226_406226 ; 
   reg __406226_406226;
   reg _406227_406227 ; 
   reg __406227_406227;
   reg _406228_406228 ; 
   reg __406228_406228;
   reg _406229_406229 ; 
   reg __406229_406229;
   reg _406230_406230 ; 
   reg __406230_406230;
   reg _406231_406231 ; 
   reg __406231_406231;
   reg _406232_406232 ; 
   reg __406232_406232;
   reg _406233_406233 ; 
   reg __406233_406233;
   reg _406234_406234 ; 
   reg __406234_406234;
   reg _406235_406235 ; 
   reg __406235_406235;
   reg _406236_406236 ; 
   reg __406236_406236;
   reg _406237_406237 ; 
   reg __406237_406237;
   reg _406238_406238 ; 
   reg __406238_406238;
   reg _406239_406239 ; 
   reg __406239_406239;
   reg _406240_406240 ; 
   reg __406240_406240;
   reg _406241_406241 ; 
   reg __406241_406241;
   reg _406242_406242 ; 
   reg __406242_406242;
   reg _406243_406243 ; 
   reg __406243_406243;
   reg _406244_406244 ; 
   reg __406244_406244;
   reg _406245_406245 ; 
   reg __406245_406245;
   reg _406246_406246 ; 
   reg __406246_406246;
   reg _406247_406247 ; 
   reg __406247_406247;
   reg _406248_406248 ; 
   reg __406248_406248;
   reg _406249_406249 ; 
   reg __406249_406249;
   reg _406250_406250 ; 
   reg __406250_406250;
   reg _406251_406251 ; 
   reg __406251_406251;
   reg _406252_406252 ; 
   reg __406252_406252;
   reg _406253_406253 ; 
   reg __406253_406253;
   reg _406254_406254 ; 
   reg __406254_406254;
   reg _406255_406255 ; 
   reg __406255_406255;
   reg _406256_406256 ; 
   reg __406256_406256;
   reg _406257_406257 ; 
   reg __406257_406257;
   reg _406258_406258 ; 
   reg __406258_406258;
   reg _406259_406259 ; 
   reg __406259_406259;
   reg _406260_406260 ; 
   reg __406260_406260;
   reg _406261_406261 ; 
   reg __406261_406261;
   reg _406262_406262 ; 
   reg __406262_406262;
   reg _406263_406263 ; 
   reg __406263_406263;
   reg _406264_406264 ; 
   reg __406264_406264;
   reg _406265_406265 ; 
   reg __406265_406265;
   reg _406266_406266 ; 
   reg __406266_406266;
   reg _406267_406267 ; 
   reg __406267_406267;
   reg _406268_406268 ; 
   reg __406268_406268;
   reg _406269_406269 ; 
   reg __406269_406269;
   reg _406270_406270 ; 
   reg __406270_406270;
   reg _406271_406271 ; 
   reg __406271_406271;
   reg _406272_406272 ; 
   reg __406272_406272;
   reg _406273_406273 ; 
   reg __406273_406273;
   reg _406274_406274 ; 
   reg __406274_406274;
   reg _406275_406275 ; 
   reg __406275_406275;
   reg _406276_406276 ; 
   reg __406276_406276;
   reg _406277_406277 ; 
   reg __406277_406277;
   reg _406278_406278 ; 
   reg __406278_406278;
   reg _406279_406279 ; 
   reg __406279_406279;
   reg _406280_406280 ; 
   reg __406280_406280;
   reg _406281_406281 ; 
   reg __406281_406281;
   reg _406282_406282 ; 
   reg __406282_406282;
   reg _406283_406283 ; 
   reg __406283_406283;
   reg _406284_406284 ; 
   reg __406284_406284;
   reg _406285_406285 ; 
   reg __406285_406285;
   reg _406286_406286 ; 
   reg __406286_406286;
   reg _406287_406287 ; 
   reg __406287_406287;
   reg _406288_406288 ; 
   reg __406288_406288;
   reg _406289_406289 ; 
   reg __406289_406289;
   reg _406290_406290 ; 
   reg __406290_406290;
   reg _406291_406291 ; 
   reg __406291_406291;
   reg _406292_406292 ; 
   reg __406292_406292;
   reg _406293_406293 ; 
   reg __406293_406293;
   reg _406294_406294 ; 
   reg __406294_406294;
   reg _406295_406295 ; 
   reg __406295_406295;
   reg _406296_406296 ; 
   reg __406296_406296;
   reg _406297_406297 ; 
   reg __406297_406297;
   reg _406298_406298 ; 
   reg __406298_406298;
   reg _406299_406299 ; 
   reg __406299_406299;
   reg _406300_406300 ; 
   reg __406300_406300;
   reg _406301_406301 ; 
   reg __406301_406301;
   reg _406302_406302 ; 
   reg __406302_406302;
   reg _406303_406303 ; 
   reg __406303_406303;
   reg _406304_406304 ; 
   reg __406304_406304;
   reg _406305_406305 ; 
   reg __406305_406305;
   reg _406306_406306 ; 
   reg __406306_406306;
   reg _406307_406307 ; 
   reg __406307_406307;
   reg _406308_406308 ; 
   reg __406308_406308;
   reg _406309_406309 ; 
   reg __406309_406309;
   reg _406310_406310 ; 
   reg __406310_406310;
   reg _406311_406311 ; 
   reg __406311_406311;
   reg _406312_406312 ; 
   reg __406312_406312;
   reg _406313_406313 ; 
   reg __406313_406313;
   reg _406314_406314 ; 
   reg __406314_406314;
   reg _406315_406315 ; 
   reg __406315_406315;
   reg _406316_406316 ; 
   reg __406316_406316;
   reg _406317_406317 ; 
   reg __406317_406317;
   reg _406318_406318 ; 
   reg __406318_406318;
   reg _406319_406319 ; 
   reg __406319_406319;
   reg _406320_406320 ; 
   reg __406320_406320;
   reg _406321_406321 ; 
   reg __406321_406321;
   reg _406322_406322 ; 
   reg __406322_406322;
   reg _406323_406323 ; 
   reg __406323_406323;
   reg _406324_406324 ; 
   reg __406324_406324;
   reg _406325_406325 ; 
   reg __406325_406325;
   reg _406326_406326 ; 
   reg __406326_406326;
   reg _406327_406327 ; 
   reg __406327_406327;
   reg _406328_406328 ; 
   reg __406328_406328;
   reg _406329_406329 ; 
   reg __406329_406329;
   reg _406330_406330 ; 
   reg __406330_406330;
   reg _406331_406331 ; 
   reg __406331_406331;
   reg _406332_406332 ; 
   reg __406332_406332;
   reg _406333_406333 ; 
   reg __406333_406333;
   reg _406334_406334 ; 
   reg __406334_406334;
   reg _406335_406335 ; 
   reg __406335_406335;
   reg _406336_406336 ; 
   reg __406336_406336;
   reg _406337_406337 ; 
   reg __406337_406337;
   reg _406338_406338 ; 
   reg __406338_406338;
   reg _406339_406339 ; 
   reg __406339_406339;
   reg _406340_406340 ; 
   reg __406340_406340;
   reg _406341_406341 ; 
   reg __406341_406341;
   reg _406342_406342 ; 
   reg __406342_406342;
   reg _406343_406343 ; 
   reg __406343_406343;
   reg _406344_406344 ; 
   reg __406344_406344;
   reg _406345_406345 ; 
   reg __406345_406345;
   reg _406346_406346 ; 
   reg __406346_406346;
   reg _406347_406347 ; 
   reg __406347_406347;
   reg _406348_406348 ; 
   reg __406348_406348;
   reg _406349_406349 ; 
   reg __406349_406349;
   reg _406350_406350 ; 
   reg __406350_406350;
   reg _406351_406351 ; 
   reg __406351_406351;
   reg _406352_406352 ; 
   reg __406352_406352;
   reg _406353_406353 ; 
   reg __406353_406353;
   reg _406354_406354 ; 
   reg __406354_406354;
   reg _406355_406355 ; 
   reg __406355_406355;
   reg _406356_406356 ; 
   reg __406356_406356;
   reg _406357_406357 ; 
   reg __406357_406357;
   reg _406358_406358 ; 
   reg __406358_406358;
   reg _406359_406359 ; 
   reg __406359_406359;
   reg _406360_406360 ; 
   reg __406360_406360;
   reg _406361_406361 ; 
   reg __406361_406361;
   reg _406362_406362 ; 
   reg __406362_406362;
   reg _406363_406363 ; 
   reg __406363_406363;
   reg _406364_406364 ; 
   reg __406364_406364;
   reg _406365_406365 ; 
   reg __406365_406365;
   reg _406366_406366 ; 
   reg __406366_406366;
   reg _406367_406367 ; 
   reg __406367_406367;
   reg _406368_406368 ; 
   reg __406368_406368;
   reg _406369_406369 ; 
   reg __406369_406369;
   reg _406370_406370 ; 
   reg __406370_406370;
   reg _406371_406371 ; 
   reg __406371_406371;
   reg _406372_406372 ; 
   reg __406372_406372;
   reg _406373_406373 ; 
   reg __406373_406373;
   reg _406374_406374 ; 
   reg __406374_406374;
   reg _406375_406375 ; 
   reg __406375_406375;
   reg _406376_406376 ; 
   reg __406376_406376;
   reg _406377_406377 ; 
   reg __406377_406377;
   reg _406378_406378 ; 
   reg __406378_406378;
   reg _406379_406379 ; 
   reg __406379_406379;
   reg _406380_406380 ; 
   reg __406380_406380;
   reg _406381_406381 ; 
   reg __406381_406381;
   reg _406382_406382 ; 
   reg __406382_406382;
   reg _406383_406383 ; 
   reg __406383_406383;
   reg _406384_406384 ; 
   reg __406384_406384;
   reg _406385_406385 ; 
   reg __406385_406385;
   reg _406386_406386 ; 
   reg __406386_406386;
   reg _406387_406387 ; 
   reg __406387_406387;
   reg _406388_406388 ; 
   reg __406388_406388;
   reg _406389_406389 ; 
   reg __406389_406389;
   reg _406390_406390 ; 
   reg __406390_406390;
   reg _406391_406391 ; 
   reg __406391_406391;
   reg _406392_406392 ; 
   reg __406392_406392;
   reg _406393_406393 ; 
   reg __406393_406393;
   reg _406394_406394 ; 
   reg __406394_406394;
   reg _406395_406395 ; 
   reg __406395_406395;
   reg _406396_406396 ; 
   reg __406396_406396;
   reg _406397_406397 ; 
   reg __406397_406397;
   reg _406398_406398 ; 
   reg __406398_406398;
   reg _406399_406399 ; 
   reg __406399_406399;
   reg _406400_406400 ; 
   reg __406400_406400;
   reg _406401_406401 ; 
   reg __406401_406401;
   reg _406402_406402 ; 
   reg __406402_406402;
   reg _406403_406403 ; 
   reg __406403_406403;
   reg _406404_406404 ; 
   reg __406404_406404;
   reg _406405_406405 ; 
   reg __406405_406405;
   reg _406406_406406 ; 
   reg __406406_406406;
   reg _406407_406407 ; 
   reg __406407_406407;
   reg _406408_406408 ; 
   reg __406408_406408;
   reg _406409_406409 ; 
   reg __406409_406409;
   reg _406410_406410 ; 
   reg __406410_406410;
   reg _406411_406411 ; 
   reg __406411_406411;
   reg _406412_406412 ; 
   reg __406412_406412;
   reg _406413_406413 ; 
   reg __406413_406413;
   reg _406414_406414 ; 
   reg __406414_406414;
   reg _406415_406415 ; 
   reg __406415_406415;
   reg _406416_406416 ; 
   reg __406416_406416;
   reg _406417_406417 ; 
   reg __406417_406417;
   reg _406418_406418 ; 
   reg __406418_406418;
   reg _406419_406419 ; 
   reg __406419_406419;
   reg _406420_406420 ; 
   reg __406420_406420;
   reg _406421_406421 ; 
   reg __406421_406421;
   reg _406422_406422 ; 
   reg __406422_406422;
   reg _406423_406423 ; 
   reg __406423_406423;
   reg _406424_406424 ; 
   reg __406424_406424;
   reg _406425_406425 ; 
   reg __406425_406425;
   reg _406426_406426 ; 
   reg __406426_406426;
   reg _406427_406427 ; 
   reg __406427_406427;
   reg _406428_406428 ; 
   reg __406428_406428;
   reg _406429_406429 ; 
   reg __406429_406429;
   reg _406430_406430 ; 
   reg __406430_406430;
   reg _406431_406431 ; 
   reg __406431_406431;
   reg _406432_406432 ; 
   reg __406432_406432;
   reg _406433_406433 ; 
   reg __406433_406433;
   reg _406434_406434 ; 
   reg __406434_406434;
   reg _406435_406435 ; 
   reg __406435_406435;
   reg _406436_406436 ; 
   reg __406436_406436;
   reg _406437_406437 ; 
   reg __406437_406437;
   reg _406438_406438 ; 
   reg __406438_406438;
   reg _406439_406439 ; 
   reg __406439_406439;
   reg _406440_406440 ; 
   reg __406440_406440;
   reg _406441_406441 ; 
   reg __406441_406441;
   reg _406442_406442 ; 
   reg __406442_406442;
   reg _406443_406443 ; 
   reg __406443_406443;
   reg _406444_406444 ; 
   reg __406444_406444;
   reg _406445_406445 ; 
   reg __406445_406445;
   reg _406446_406446 ; 
   reg __406446_406446;
   reg _406447_406447 ; 
   reg __406447_406447;
   reg _406448_406448 ; 
   reg __406448_406448;
   reg _406449_406449 ; 
   reg __406449_406449;
   reg _406450_406450 ; 
   reg __406450_406450;
   reg _406451_406451 ; 
   reg __406451_406451;
   reg _406452_406452 ; 
   reg __406452_406452;
   reg _406453_406453 ; 
   reg __406453_406453;
   reg _406454_406454 ; 
   reg __406454_406454;
   reg _406455_406455 ; 
   reg __406455_406455;
   reg _406456_406456 ; 
   reg __406456_406456;
   reg _406457_406457 ; 
   reg __406457_406457;
   reg _406458_406458 ; 
   reg __406458_406458;
   reg _406459_406459 ; 
   reg __406459_406459;
   reg _406460_406460 ; 
   reg __406460_406460;
   reg _406461_406461 ; 
   reg __406461_406461;
   reg _406462_406462 ; 
   reg __406462_406462;
   reg _406463_406463 ; 
   reg __406463_406463;
   reg _406464_406464 ; 
   reg __406464_406464;
   reg _406465_406465 ; 
   reg __406465_406465;
   reg _406466_406466 ; 
   reg __406466_406466;
   reg _406467_406467 ; 
   reg __406467_406467;
   reg _406468_406468 ; 
   reg __406468_406468;
   reg _406469_406469 ; 
   reg __406469_406469;
   reg _406470_406470 ; 
   reg __406470_406470;
   reg _406471_406471 ; 
   reg __406471_406471;
   reg _406472_406472 ; 
   reg __406472_406472;
   reg _406473_406473 ; 
   reg __406473_406473;
   reg _406474_406474 ; 
   reg __406474_406474;
   reg _406475_406475 ; 
   reg __406475_406475;
   reg _406476_406476 ; 
   reg __406476_406476;
   reg _406477_406477 ; 
   reg __406477_406477;
   reg _406478_406478 ; 
   reg __406478_406478;
   reg _406479_406479 ; 
   reg __406479_406479;
   reg _406480_406480 ; 
   reg __406480_406480;
   reg _406481_406481 ; 
   reg __406481_406481;
   reg _406482_406482 ; 
   reg __406482_406482;
   reg _406483_406483 ; 
   reg __406483_406483;
   reg _406484_406484 ; 
   reg __406484_406484;
   reg _406485_406485 ; 
   reg __406485_406485;
   reg _406486_406486 ; 
   reg __406486_406486;
   reg _406487_406487 ; 
   reg __406487_406487;
   reg _406488_406488 ; 
   reg __406488_406488;
   reg _406489_406489 ; 
   reg __406489_406489;
   reg _406490_406490 ; 
   reg __406490_406490;
   reg _406491_406491 ; 
   reg __406491_406491;
   reg _406492_406492 ; 
   reg __406492_406492;
   reg _406493_406493 ; 
   reg __406493_406493;
   reg _406494_406494 ; 
   reg __406494_406494;
   reg _406495_406495 ; 
   reg __406495_406495;
   reg _406496_406496 ; 
   reg __406496_406496;
   reg _406497_406497 ; 
   reg __406497_406497;
   reg _406498_406498 ; 
   reg __406498_406498;
   reg _406499_406499 ; 
   reg __406499_406499;
   reg _406500_406500 ; 
   reg __406500_406500;
   reg _406501_406501 ; 
   reg __406501_406501;
   reg _406502_406502 ; 
   reg __406502_406502;
   reg _406503_406503 ; 
   reg __406503_406503;
   reg _406504_406504 ; 
   reg __406504_406504;
   reg _406505_406505 ; 
   reg __406505_406505;
   reg _406506_406506 ; 
   reg __406506_406506;
   reg _406507_406507 ; 
   reg __406507_406507;
   reg _406508_406508 ; 
   reg __406508_406508;
   reg _406509_406509 ; 
   reg __406509_406509;
   reg _406510_406510 ; 
   reg __406510_406510;
   reg _406511_406511 ; 
   reg __406511_406511;
   reg _406512_406512 ; 
   reg __406512_406512;
   reg _406513_406513 ; 
   reg __406513_406513;
   reg _406514_406514 ; 
   reg __406514_406514;
   reg _406515_406515 ; 
   reg __406515_406515;
   reg _406516_406516 ; 
   reg __406516_406516;
   reg _406517_406517 ; 
   reg __406517_406517;
   reg _406518_406518 ; 
   reg __406518_406518;
   reg _406519_406519 ; 
   reg __406519_406519;
   reg _406520_406520 ; 
   reg __406520_406520;
   reg _406521_406521 ; 
   reg __406521_406521;
   reg _406522_406522 ; 
   reg __406522_406522;
   reg _406523_406523 ; 
   reg __406523_406523;
   reg _406524_406524 ; 
   reg __406524_406524;
   reg _406525_406525 ; 
   reg __406525_406525;
   reg _406526_406526 ; 
   reg __406526_406526;
   reg _406527_406527 ; 
   reg __406527_406527;
   reg _406528_406528 ; 
   reg __406528_406528;
   reg _406529_406529 ; 
   reg __406529_406529;
   reg _406530_406530 ; 
   reg __406530_406530;
   reg _406531_406531 ; 
   reg __406531_406531;
   reg _406532_406532 ; 
   reg __406532_406532;
   reg _406533_406533 ; 
   reg __406533_406533;
   reg _406534_406534 ; 
   reg __406534_406534;
   reg _406535_406535 ; 
   reg __406535_406535;
   reg _406536_406536 ; 
   reg __406536_406536;
   reg _406537_406537 ; 
   reg __406537_406537;
   reg _406538_406538 ; 
   reg __406538_406538;
   reg _406539_406539 ; 
   reg __406539_406539;
   reg _406540_406540 ; 
   reg __406540_406540;
   reg _406541_406541 ; 
   reg __406541_406541;
   reg _406542_406542 ; 
   reg __406542_406542;
   reg _406543_406543 ; 
   reg __406543_406543;
   reg _406544_406544 ; 
   reg __406544_406544;
   reg _406545_406545 ; 
   reg __406545_406545;
   reg _406546_406546 ; 
   reg __406546_406546;
   reg _406547_406547 ; 
   reg __406547_406547;
   reg _406548_406548 ; 
   reg __406548_406548;
   reg _406549_406549 ; 
   reg __406549_406549;
   reg _406550_406550 ; 
   reg __406550_406550;
   reg _406551_406551 ; 
   reg __406551_406551;
   reg _406552_406552 ; 
   reg __406552_406552;
   reg _406553_406553 ; 
   reg __406553_406553;
   reg _406554_406554 ; 
   reg __406554_406554;
   reg _406555_406555 ; 
   reg __406555_406555;
   reg _406556_406556 ; 
   reg __406556_406556;
   reg _406557_406557 ; 
   reg __406557_406557;
   reg _406558_406558 ; 
   reg __406558_406558;
   reg _406559_406559 ; 
   reg __406559_406559;
   reg _406560_406560 ; 
   reg __406560_406560;
   reg _406561_406561 ; 
   reg __406561_406561;
   reg _406562_406562 ; 
   reg __406562_406562;
   reg _406563_406563 ; 
   reg __406563_406563;
   reg _406564_406564 ; 
   reg __406564_406564;
   reg _406565_406565 ; 
   reg __406565_406565;
   reg _406566_406566 ; 
   reg __406566_406566;
   reg _406567_406567 ; 
   reg __406567_406567;
   reg _406568_406568 ; 
   reg __406568_406568;
   reg _406569_406569 ; 
   reg __406569_406569;
   reg _406570_406570 ; 
   reg __406570_406570;
   reg _406571_406571 ; 
   reg __406571_406571;
   reg _406572_406572 ; 
   reg __406572_406572;
   reg _406573_406573 ; 
   reg __406573_406573;
   reg _406574_406574 ; 
   reg __406574_406574;
   reg _406575_406575 ; 
   reg __406575_406575;
   reg _406576_406576 ; 
   reg __406576_406576;
   reg _406577_406577 ; 
   reg __406577_406577;
   reg _406578_406578 ; 
   reg __406578_406578;
   reg _406579_406579 ; 
   reg __406579_406579;
   reg _406580_406580 ; 
   reg __406580_406580;
   reg _406581_406581 ; 
   reg __406581_406581;
   reg _406582_406582 ; 
   reg __406582_406582;
   reg _406583_406583 ; 
   reg __406583_406583;
   reg _406584_406584 ; 
   reg __406584_406584;
   reg _406585_406585 ; 
   reg __406585_406585;
   reg _406586_406586 ; 
   reg __406586_406586;
   reg _406587_406587 ; 
   reg __406587_406587;
   reg _406588_406588 ; 
   reg __406588_406588;
   reg _406589_406589 ; 
   reg __406589_406589;
   reg _406590_406590 ; 
   reg __406590_406590;
   reg _406591_406591 ; 
   reg __406591_406591;
   reg _406592_406592 ; 
   reg __406592_406592;
   reg _406593_406593 ; 
   reg __406593_406593;
   reg _406594_406594 ; 
   reg __406594_406594;
   reg _406595_406595 ; 
   reg __406595_406595;
   reg _406596_406596 ; 
   reg __406596_406596;
   reg _406597_406597 ; 
   reg __406597_406597;
   reg _406598_406598 ; 
   reg __406598_406598;
   reg _406599_406599 ; 
   reg __406599_406599;
   reg _406600_406600 ; 
   reg __406600_406600;
   reg _406601_406601 ; 
   reg __406601_406601;
   reg _406602_406602 ; 
   reg __406602_406602;
   reg _406603_406603 ; 
   reg __406603_406603;
   reg _406604_406604 ; 
   reg __406604_406604;
   reg _406605_406605 ; 
   reg __406605_406605;
   reg _406606_406606 ; 
   reg __406606_406606;
   reg _406607_406607 ; 
   reg __406607_406607;
   reg _406608_406608 ; 
   reg __406608_406608;
   reg _406609_406609 ; 
   reg __406609_406609;
   reg _406610_406610 ; 
   reg __406610_406610;
   reg _406611_406611 ; 
   reg __406611_406611;
   reg _406612_406612 ; 
   reg __406612_406612;
   reg _406613_406613 ; 
   reg __406613_406613;
   reg _406614_406614 ; 
   reg __406614_406614;
   reg _406615_406615 ; 
   reg __406615_406615;
   reg _406616_406616 ; 
   reg __406616_406616;
   reg _406617_406617 ; 
   reg __406617_406617;
   reg _406618_406618 ; 
   reg __406618_406618;
   reg _406619_406619 ; 
   reg __406619_406619;
   reg _406620_406620 ; 
   reg __406620_406620;
   reg _406621_406621 ; 
   reg __406621_406621;
   reg _406622_406622 ; 
   reg __406622_406622;
   reg _406623_406623 ; 
   reg __406623_406623;
   reg _406624_406624 ; 
   reg __406624_406624;
   reg _406625_406625 ; 
   reg __406625_406625;
   reg _406626_406626 ; 
   reg __406626_406626;
   reg _406627_406627 ; 
   reg __406627_406627;
   reg _406628_406628 ; 
   reg __406628_406628;
   reg _406629_406629 ; 
   reg __406629_406629;
   reg _406630_406630 ; 
   reg __406630_406630;
   reg _406631_406631 ; 
   reg __406631_406631;
   reg _406632_406632 ; 
   reg __406632_406632;
   reg _406633_406633 ; 
   reg __406633_406633;
   reg _406634_406634 ; 
   reg __406634_406634;
   reg _406635_406635 ; 
   reg __406635_406635;
   reg _406636_406636 ; 
   reg __406636_406636;
   reg _406637_406637 ; 
   reg __406637_406637;
   reg _406638_406638 ; 
   reg __406638_406638;
   reg _406639_406639 ; 
   reg __406639_406639;
   reg _406640_406640 ; 
   reg __406640_406640;
   reg _406641_406641 ; 
   reg __406641_406641;
   reg _406642_406642 ; 
   reg __406642_406642;
   reg _406643_406643 ; 
   reg __406643_406643;
   reg _406644_406644 ; 
   reg __406644_406644;
   reg _406645_406645 ; 
   reg __406645_406645;
   reg _406646_406646 ; 
   reg __406646_406646;
   reg _406647_406647 ; 
   reg __406647_406647;
   reg _406648_406648 ; 
   reg __406648_406648;
   reg _406649_406649 ; 
   reg __406649_406649;
   reg _406650_406650 ; 
   reg __406650_406650;
   reg _406651_406651 ; 
   reg __406651_406651;
   reg _406652_406652 ; 
   reg __406652_406652;
   reg _406653_406653 ; 
   reg __406653_406653;
   reg _406654_406654 ; 
   reg __406654_406654;
   reg _406655_406655 ; 
   reg __406655_406655;
   reg _406656_406656 ; 
   reg __406656_406656;
   reg _406657_406657 ; 
   reg __406657_406657;
   reg _406658_406658 ; 
   reg __406658_406658;
   reg _406659_406659 ; 
   reg __406659_406659;
   reg _406660_406660 ; 
   reg __406660_406660;
   reg _406661_406661 ; 
   reg __406661_406661;
   reg _406662_406662 ; 
   reg __406662_406662;
   reg _406663_406663 ; 
   reg __406663_406663;
   reg _406664_406664 ; 
   reg __406664_406664;
   reg _406665_406665 ; 
   reg __406665_406665;
   reg _406666_406666 ; 
   reg __406666_406666;
   reg _406667_406667 ; 
   reg __406667_406667;
   reg _406668_406668 ; 
   reg __406668_406668;
   reg _406669_406669 ; 
   reg __406669_406669;
   reg _406670_406670 ; 
   reg __406670_406670;
   reg _406671_406671 ; 
   reg __406671_406671;
   reg _406672_406672 ; 
   reg __406672_406672;
   reg _406673_406673 ; 
   reg __406673_406673;
   reg _406674_406674 ; 
   reg __406674_406674;
   reg _406675_406675 ; 
   reg __406675_406675;
   reg _406676_406676 ; 
   reg __406676_406676;
   reg _406677_406677 ; 
   reg __406677_406677;
   reg _406678_406678 ; 
   reg __406678_406678;
   reg _406679_406679 ; 
   reg __406679_406679;
   reg _406680_406680 ; 
   reg __406680_406680;
   reg _406681_406681 ; 
   reg __406681_406681;
   reg _406682_406682 ; 
   reg __406682_406682;
   reg _406683_406683 ; 
   reg __406683_406683;
   reg _406684_406684 ; 
   reg __406684_406684;
   reg _406685_406685 ; 
   reg __406685_406685;
   reg _406686_406686 ; 
   reg __406686_406686;
   reg _406687_406687 ; 
   reg __406687_406687;
   reg _406688_406688 ; 
   reg __406688_406688;
   reg _406689_406689 ; 
   reg __406689_406689;
   reg _406690_406690 ; 
   reg __406690_406690;
   reg _406691_406691 ; 
   reg __406691_406691;
   reg _406692_406692 ; 
   reg __406692_406692;
   reg _406693_406693 ; 
   reg __406693_406693;
   reg _406694_406694 ; 
   reg __406694_406694;
   reg _406695_406695 ; 
   reg __406695_406695;
   reg _406696_406696 ; 
   reg __406696_406696;
   reg _406697_406697 ; 
   reg __406697_406697;
   reg _406698_406698 ; 
   reg __406698_406698;
   reg _406699_406699 ; 
   reg __406699_406699;
   reg _406700_406700 ; 
   reg __406700_406700;
   reg _406701_406701 ; 
   reg __406701_406701;
   reg _406702_406702 ; 
   reg __406702_406702;
   reg _406703_406703 ; 
   reg __406703_406703;
   reg _406704_406704 ; 
   reg __406704_406704;
   reg _406705_406705 ; 
   reg __406705_406705;
   reg _406706_406706 ; 
   reg __406706_406706;
   reg _406707_406707 ; 
   reg __406707_406707;
   reg _406708_406708 ; 
   reg __406708_406708;
   reg _406709_406709 ; 
   reg __406709_406709;
   reg _406710_406710 ; 
   reg __406710_406710;
   reg _406711_406711 ; 
   reg __406711_406711;
   reg _406712_406712 ; 
   reg __406712_406712;
   reg _406713_406713 ; 
   reg __406713_406713;
   reg _406714_406714 ; 
   reg __406714_406714;
   reg _406715_406715 ; 
   reg __406715_406715;
   reg _406716_406716 ; 
   reg __406716_406716;
   reg _406717_406717 ; 
   reg __406717_406717;
   reg _406718_406718 ; 
   reg __406718_406718;
   reg _406719_406719 ; 
   reg __406719_406719;
   reg _406720_406720 ; 
   reg __406720_406720;
   reg _406721_406721 ; 
   reg __406721_406721;
   reg _406722_406722 ; 
   reg __406722_406722;
   reg _406723_406723 ; 
   reg __406723_406723;
   reg _406724_406724 ; 
   reg __406724_406724;
   reg _406725_406725 ; 
   reg __406725_406725;
   reg _406726_406726 ; 
   reg __406726_406726;
   reg _406727_406727 ; 
   reg __406727_406727;
   reg _406728_406728 ; 
   reg __406728_406728;
   reg _406729_406729 ; 
   reg __406729_406729;
   reg _406730_406730 ; 
   reg __406730_406730;
   reg _406731_406731 ; 
   reg __406731_406731;
   reg _406732_406732 ; 
   reg __406732_406732;
   reg _406733_406733 ; 
   reg __406733_406733;
   reg _406734_406734 ; 
   reg __406734_406734;
   reg _406735_406735 ; 
   reg __406735_406735;
   reg _406736_406736 ; 
   reg __406736_406736;
   reg _406737_406737 ; 
   reg __406737_406737;
   reg _406738_406738 ; 
   reg __406738_406738;
   reg _406739_406739 ; 
   reg __406739_406739;
   reg _406740_406740 ; 
   reg __406740_406740;
   reg _406741_406741 ; 
   reg __406741_406741;
   reg _406742_406742 ; 
   reg __406742_406742;
   reg _406743_406743 ; 
   reg __406743_406743;
   reg _406744_406744 ; 
   reg __406744_406744;
   reg _406745_406745 ; 
   reg __406745_406745;
   reg _406746_406746 ; 
   reg __406746_406746;
   reg _406747_406747 ; 
   reg __406747_406747;
   reg _406748_406748 ; 
   reg __406748_406748;
   reg _406749_406749 ; 
   reg __406749_406749;
   reg _406750_406750 ; 
   reg __406750_406750;
   reg _406751_406751 ; 
   reg __406751_406751;
   reg _406752_406752 ; 
   reg __406752_406752;
   reg _406753_406753 ; 
   reg __406753_406753;
   reg _406754_406754 ; 
   reg __406754_406754;
   reg _406755_406755 ; 
   reg __406755_406755;
   reg _406756_406756 ; 
   reg __406756_406756;
   reg _406757_406757 ; 
   reg __406757_406757;
   reg _406758_406758 ; 
   reg __406758_406758;
   reg _406759_406759 ; 
   reg __406759_406759;
   reg _406760_406760 ; 
   reg __406760_406760;
   reg _406761_406761 ; 
   reg __406761_406761;
   reg _406762_406762 ; 
   reg __406762_406762;
   reg _406763_406763 ; 
   reg __406763_406763;
   reg _406764_406764 ; 
   reg __406764_406764;
   reg _406765_406765 ; 
   reg __406765_406765;
   reg _406766_406766 ; 
   reg __406766_406766;
   reg _406767_406767 ; 
   reg __406767_406767;
   reg _406768_406768 ; 
   reg __406768_406768;
   reg _406769_406769 ; 
   reg __406769_406769;
   reg _406770_406770 ; 
   reg __406770_406770;
   reg _406771_406771 ; 
   reg __406771_406771;
   reg _406772_406772 ; 
   reg __406772_406772;
   reg _406773_406773 ; 
   reg __406773_406773;
   reg _406774_406774 ; 
   reg __406774_406774;
   reg _406775_406775 ; 
   reg __406775_406775;
   reg _406776_406776 ; 
   reg __406776_406776;
   reg _406777_406777 ; 
   reg __406777_406777;
   reg _406778_406778 ; 
   reg __406778_406778;
   reg _406779_406779 ; 
   reg __406779_406779;
   reg _406780_406780 ; 
   reg __406780_406780;
   reg _406781_406781 ; 
   reg __406781_406781;
   reg _406782_406782 ; 
   reg __406782_406782;
   reg _406783_406783 ; 
   reg __406783_406783;
   reg _406784_406784 ; 
   reg __406784_406784;
   reg _406785_406785 ; 
   reg __406785_406785;
   reg _406786_406786 ; 
   reg __406786_406786;
   reg _406787_406787 ; 
   reg __406787_406787;
   reg _406788_406788 ; 
   reg __406788_406788;
   reg _406789_406789 ; 
   reg __406789_406789;
   reg _406790_406790 ; 
   reg __406790_406790;
   reg _406791_406791 ; 
   reg __406791_406791;
   reg _406792_406792 ; 
   reg __406792_406792;
   reg _406793_406793 ; 
   reg __406793_406793;
   reg _406794_406794 ; 
   reg __406794_406794;
   reg _406795_406795 ; 
   reg __406795_406795;
   reg _406796_406796 ; 
   reg __406796_406796;
   reg _406797_406797 ; 
   reg __406797_406797;
   reg _406798_406798 ; 
   reg __406798_406798;
   reg _406799_406799 ; 
   reg __406799_406799;
   reg _406800_406800 ; 
   reg __406800_406800;
   reg _406801_406801 ; 
   reg __406801_406801;
   reg _406802_406802 ; 
   reg __406802_406802;
   reg _406803_406803 ; 
   reg __406803_406803;
   reg _406804_406804 ; 
   reg __406804_406804;
   reg _406805_406805 ; 
   reg __406805_406805;
   reg _406806_406806 ; 
   reg __406806_406806;
   reg _406807_406807 ; 
   reg __406807_406807;
   reg _406808_406808 ; 
   reg __406808_406808;
   reg _406809_406809 ; 
   reg __406809_406809;
   reg _406810_406810 ; 
   reg __406810_406810;
   reg _406811_406811 ; 
   reg __406811_406811;
   reg _406812_406812 ; 
   reg __406812_406812;
   reg _406813_406813 ; 
   reg __406813_406813;
   reg _406814_406814 ; 
   reg __406814_406814;
   reg _406815_406815 ; 
   reg __406815_406815;
   reg _406816_406816 ; 
   reg __406816_406816;
   reg _406817_406817 ; 
   reg __406817_406817;
   reg _406818_406818 ; 
   reg __406818_406818;
   reg _406819_406819 ; 
   reg __406819_406819;
   reg _406820_406820 ; 
   reg __406820_406820;
   reg _406821_406821 ; 
   reg __406821_406821;
   reg _406822_406822 ; 
   reg __406822_406822;
   reg _406823_406823 ; 
   reg __406823_406823;
   reg _406824_406824 ; 
   reg __406824_406824;
   reg _406825_406825 ; 
   reg __406825_406825;
   reg _406826_406826 ; 
   reg __406826_406826;
   reg _406827_406827 ; 
   reg __406827_406827;
   reg _406828_406828 ; 
   reg __406828_406828;
   reg _406829_406829 ; 
   reg __406829_406829;
   reg _406830_406830 ; 
   reg __406830_406830;
   reg _406831_406831 ; 
   reg __406831_406831;
   reg _406832_406832 ; 
   reg __406832_406832;
   reg _406833_406833 ; 
   reg __406833_406833;
   reg _406834_406834 ; 
   reg __406834_406834;
   reg _406835_406835 ; 
   reg __406835_406835;
   reg _406836_406836 ; 
   reg __406836_406836;
   reg _406837_406837 ; 
   reg __406837_406837;
   reg _406838_406838 ; 
   reg __406838_406838;
   reg _406839_406839 ; 
   reg __406839_406839;
   reg _406840_406840 ; 
   reg __406840_406840;
   reg _406841_406841 ; 
   reg __406841_406841;
   reg _406842_406842 ; 
   reg __406842_406842;
   reg _406843_406843 ; 
   reg __406843_406843;
   reg _406844_406844 ; 
   reg __406844_406844;
   reg _406845_406845 ; 
   reg __406845_406845;
   reg _406846_406846 ; 
   reg __406846_406846;
   reg _406847_406847 ; 
   reg __406847_406847;
   reg _406848_406848 ; 
   reg __406848_406848;
   reg _406849_406849 ; 
   reg __406849_406849;
   reg _406850_406850 ; 
   reg __406850_406850;
   reg _406851_406851 ; 
   reg __406851_406851;
   reg _406852_406852 ; 
   reg __406852_406852;
   reg _406853_406853 ; 
   reg __406853_406853;
   reg _406854_406854 ; 
   reg __406854_406854;
   reg _406855_406855 ; 
   reg __406855_406855;
   reg _406856_406856 ; 
   reg __406856_406856;
   reg _406857_406857 ; 
   reg __406857_406857;
   reg _406858_406858 ; 
   reg __406858_406858;
   reg _406859_406859 ; 
   reg __406859_406859;
   reg _406860_406860 ; 
   reg __406860_406860;
   reg _406861_406861 ; 
   reg __406861_406861;
   reg _406862_406862 ; 
   reg __406862_406862;
   reg _406863_406863 ; 
   reg __406863_406863;
   reg _406864_406864 ; 
   reg __406864_406864;
   reg _406865_406865 ; 
   reg __406865_406865;
   reg _406866_406866 ; 
   reg __406866_406866;
   reg _406867_406867 ; 
   reg __406867_406867;
   reg _406868_406868 ; 
   reg __406868_406868;
   reg _406869_406869 ; 
   reg __406869_406869;
   reg _406870_406870 ; 
   reg __406870_406870;
   reg _406871_406871 ; 
   reg __406871_406871;
   reg _406872_406872 ; 
   reg __406872_406872;
   reg _406873_406873 ; 
   reg __406873_406873;
   reg _406874_406874 ; 
   reg __406874_406874;
   reg _406875_406875 ; 
   reg __406875_406875;
   reg _406876_406876 ; 
   reg __406876_406876;
   reg _406877_406877 ; 
   reg __406877_406877;
   reg _406878_406878 ; 
   reg __406878_406878;
   reg _406879_406879 ; 
   reg __406879_406879;
   reg _406880_406880 ; 
   reg __406880_406880;
   reg _406881_406881 ; 
   reg __406881_406881;
   reg _406882_406882 ; 
   reg __406882_406882;
   reg _406883_406883 ; 
   reg __406883_406883;
   reg _406884_406884 ; 
   reg __406884_406884;
   reg _406885_406885 ; 
   reg __406885_406885;
   reg _406886_406886 ; 
   reg __406886_406886;
   reg _406887_406887 ; 
   reg __406887_406887;
   reg _406888_406888 ; 
   reg __406888_406888;
   reg _406889_406889 ; 
   reg __406889_406889;
   reg _406890_406890 ; 
   reg __406890_406890;
   reg _406891_406891 ; 
   reg __406891_406891;
   reg _406892_406892 ; 
   reg __406892_406892;
   reg _406893_406893 ; 
   reg __406893_406893;
   reg _406894_406894 ; 
   reg __406894_406894;
   reg _406895_406895 ; 
   reg __406895_406895;
   reg _406896_406896 ; 
   reg __406896_406896;
   reg _406897_406897 ; 
   reg __406897_406897;
   reg _406898_406898 ; 
   reg __406898_406898;
   reg _406899_406899 ; 
   reg __406899_406899;
   reg _406900_406900 ; 
   reg __406900_406900;
   reg _406901_406901 ; 
   reg __406901_406901;
   reg _406902_406902 ; 
   reg __406902_406902;
   reg _406903_406903 ; 
   reg __406903_406903;
   reg _406904_406904 ; 
   reg __406904_406904;
   reg _406905_406905 ; 
   reg __406905_406905;
   reg _406906_406906 ; 
   reg __406906_406906;
   reg _406907_406907 ; 
   reg __406907_406907;
   reg _406908_406908 ; 
   reg __406908_406908;
   reg _406909_406909 ; 
   reg __406909_406909;
   reg _406910_406910 ; 
   reg __406910_406910;
   reg _406911_406911 ; 
   reg __406911_406911;
   reg _406912_406912 ; 
   reg __406912_406912;
   reg _406913_406913 ; 
   reg __406913_406913;
   reg _406914_406914 ; 
   reg __406914_406914;
   reg _406915_406915 ; 
   reg __406915_406915;
   reg _406916_406916 ; 
   reg __406916_406916;
   reg _406917_406917 ; 
   reg __406917_406917;
   reg _406918_406918 ; 
   reg __406918_406918;
   reg _406919_406919 ; 
   reg __406919_406919;
   reg _406920_406920 ; 
   reg __406920_406920;
   reg _406921_406921 ; 
   reg __406921_406921;
   reg _406922_406922 ; 
   reg __406922_406922;
   reg _406923_406923 ; 
   reg __406923_406923;
   reg _406924_406924 ; 
   reg __406924_406924;
   reg _406925_406925 ; 
   reg __406925_406925;
   reg _406926_406926 ; 
   reg __406926_406926;
   reg _406927_406927 ; 
   reg __406927_406927;
   reg _406928_406928 ; 
   reg __406928_406928;
   reg _406929_406929 ; 
   reg __406929_406929;
   reg _406930_406930 ; 
   reg __406930_406930;
   reg _406931_406931 ; 
   reg __406931_406931;
   reg _406932_406932 ; 
   reg __406932_406932;
   reg _406933_406933 ; 
   reg __406933_406933;
   reg _406934_406934 ; 
   reg __406934_406934;
   reg _406935_406935 ; 
   reg __406935_406935;
   reg _406936_406936 ; 
   reg __406936_406936;
   reg _406937_406937 ; 
   reg __406937_406937;
   reg _406938_406938 ; 
   reg __406938_406938;
   reg _406939_406939 ; 
   reg __406939_406939;
   reg _406940_406940 ; 
   reg __406940_406940;
   reg _406941_406941 ; 
   reg __406941_406941;
   reg _406942_406942 ; 
   reg __406942_406942;
   reg _406943_406943 ; 
   reg __406943_406943;
   reg _406944_406944 ; 
   reg __406944_406944;
   reg _406945_406945 ; 
   reg __406945_406945;
   reg _406946_406946 ; 
   reg __406946_406946;
   reg _406947_406947 ; 
   reg __406947_406947;
   reg _406948_406948 ; 
   reg __406948_406948;
   reg _406949_406949 ; 
   reg __406949_406949;
   reg _406950_406950 ; 
   reg __406950_406950;
   reg _406951_406951 ; 
   reg __406951_406951;
   reg _406952_406952 ; 
   reg __406952_406952;
   reg _406953_406953 ; 
   reg __406953_406953;
   reg _406954_406954 ; 
   reg __406954_406954;
   reg _406955_406955 ; 
   reg __406955_406955;
   reg _406956_406956 ; 
   reg __406956_406956;
   reg _406957_406957 ; 
   reg __406957_406957;
   reg _406958_406958 ; 
   reg __406958_406958;
   reg _406959_406959 ; 
   reg __406959_406959;
   reg _406960_406960 ; 
   reg __406960_406960;
   reg _406961_406961 ; 
   reg __406961_406961;
   reg _406962_406962 ; 
   reg __406962_406962;
   reg _406963_406963 ; 
   reg __406963_406963;
   reg _406964_406964 ; 
   reg __406964_406964;
   reg _406965_406965 ; 
   reg __406965_406965;
   reg _406966_406966 ; 
   reg __406966_406966;
   reg _406967_406967 ; 
   reg __406967_406967;
   reg _406968_406968 ; 
   reg __406968_406968;
   reg _406969_406969 ; 
   reg __406969_406969;
   reg _406970_406970 ; 
   reg __406970_406970;
   reg _406971_406971 ; 
   reg __406971_406971;
   reg _406972_406972 ; 
   reg __406972_406972;
   reg _406973_406973 ; 
   reg __406973_406973;
   reg _406974_406974 ; 
   reg __406974_406974;
   reg _406975_406975 ; 
   reg __406975_406975;
   reg _406976_406976 ; 
   reg __406976_406976;
   reg _406977_406977 ; 
   reg __406977_406977;
   reg _406978_406978 ; 
   reg __406978_406978;
   reg _406979_406979 ; 
   reg __406979_406979;
   reg _406980_406980 ; 
   reg __406980_406980;
   reg _406981_406981 ; 
   reg __406981_406981;
   reg _406982_406982 ; 
   reg __406982_406982;
   reg _406983_406983 ; 
   reg __406983_406983;
   reg _406984_406984 ; 
   reg __406984_406984;
   reg _406985_406985 ; 
   reg __406985_406985;
   reg _406986_406986 ; 
   reg __406986_406986;
   reg _406987_406987 ; 
   reg __406987_406987;
   reg _406988_406988 ; 
   reg __406988_406988;
   reg _406989_406989 ; 
   reg __406989_406989;
   reg _406990_406990 ; 
   reg __406990_406990;
   reg _406991_406991 ; 
   reg __406991_406991;
   reg _406992_406992 ; 
   reg __406992_406992;
   reg _406993_406993 ; 
   reg __406993_406993;
   reg _406994_406994 ; 
   reg __406994_406994;
   reg _406995_406995 ; 
   reg __406995_406995;
   reg _406996_406996 ; 
   reg __406996_406996;
   reg _406997_406997 ; 
   reg __406997_406997;
   reg _406998_406998 ; 
   reg __406998_406998;
   reg _406999_406999 ; 
   reg __406999_406999;
   reg _407000_407000 ; 
   reg __407000_407000;
   reg _407001_407001 ; 
   reg __407001_407001;
   reg _407002_407002 ; 
   reg __407002_407002;
   reg _407003_407003 ; 
   reg __407003_407003;
   reg _407004_407004 ; 
   reg __407004_407004;
   reg _407005_407005 ; 
   reg __407005_407005;
   reg _407006_407006 ; 
   reg __407006_407006;
   reg _407007_407007 ; 
   reg __407007_407007;
   reg _407008_407008 ; 
   reg __407008_407008;
   reg _407009_407009 ; 
   reg __407009_407009;
   reg _407010_407010 ; 
   reg __407010_407010;
   reg _407011_407011 ; 
   reg __407011_407011;
   reg _407012_407012 ; 
   reg __407012_407012;
   reg _407013_407013 ; 
   reg __407013_407013;
   reg _407014_407014 ; 
   reg __407014_407014;
   reg _407015_407015 ; 
   reg __407015_407015;
   reg _407016_407016 ; 
   reg __407016_407016;
   reg _407017_407017 ; 
   reg __407017_407017;
   reg _407018_407018 ; 
   reg __407018_407018;
   reg _407019_407019 ; 
   reg __407019_407019;
   reg _407020_407020 ; 
   reg __407020_407020;
   reg _407021_407021 ; 
   reg __407021_407021;
   reg _407022_407022 ; 
   reg __407022_407022;
   reg _407023_407023 ; 
   reg __407023_407023;
   reg _407024_407024 ; 
   reg __407024_407024;
   reg _407025_407025 ; 
   reg __407025_407025;
   reg _407026_407026 ; 
   reg __407026_407026;
   reg _407027_407027 ; 
   reg __407027_407027;
   reg _407028_407028 ; 
   reg __407028_407028;
   reg _407029_407029 ; 
   reg __407029_407029;
   reg _407030_407030 ; 
   reg __407030_407030;
   reg _407031_407031 ; 
   reg __407031_407031;
   reg _407032_407032 ; 
   reg __407032_407032;
   reg _407033_407033 ; 
   reg __407033_407033;
   reg _407034_407034 ; 
   reg __407034_407034;
   reg _407035_407035 ; 
   reg __407035_407035;
   reg _407036_407036 ; 
   reg __407036_407036;
   reg _407037_407037 ; 
   reg __407037_407037;
   reg _407038_407038 ; 
   reg __407038_407038;
   reg _407039_407039 ; 
   reg __407039_407039;
   reg _407040_407040 ; 
   reg __407040_407040;
   reg _407041_407041 ; 
   reg __407041_407041;
   reg _407042_407042 ; 
   reg __407042_407042;
   reg _407043_407043 ; 
   reg __407043_407043;
   reg _407044_407044 ; 
   reg __407044_407044;
   reg _407045_407045 ; 
   reg __407045_407045;
   reg _407046_407046 ; 
   reg __407046_407046;
   reg _407047_407047 ; 
   reg __407047_407047;
   reg _407048_407048 ; 
   reg __407048_407048;
   reg _407049_407049 ; 
   reg __407049_407049;
   reg _407050_407050 ; 
   reg __407050_407050;
   reg _407051_407051 ; 
   reg __407051_407051;
   reg _407052_407052 ; 
   reg __407052_407052;
   reg _407053_407053 ; 
   reg __407053_407053;
   reg _407054_407054 ; 
   reg __407054_407054;
   reg _407055_407055 ; 
   reg __407055_407055;
   reg _407056_407056 ; 
   reg __407056_407056;
   reg _407057_407057 ; 
   reg __407057_407057;
   reg _407058_407058 ; 
   reg __407058_407058;
   reg _407059_407059 ; 
   reg __407059_407059;
   reg _407060_407060 ; 
   reg __407060_407060;
   reg _407061_407061 ; 
   reg __407061_407061;
   reg _407062_407062 ; 
   reg __407062_407062;
   reg _407063_407063 ; 
   reg __407063_407063;
   reg _407064_407064 ; 
   reg __407064_407064;
   reg _407065_407065 ; 
   reg __407065_407065;
   reg _407066_407066 ; 
   reg __407066_407066;
   reg _407067_407067 ; 
   reg __407067_407067;
   reg _407068_407068 ; 
   reg __407068_407068;
   reg _407069_407069 ; 
   reg __407069_407069;
   reg _407070_407070 ; 
   reg __407070_407070;
   reg _407071_407071 ; 
   reg __407071_407071;
   reg _407072_407072 ; 
   reg __407072_407072;
   reg _407073_407073 ; 
   reg __407073_407073;
   reg _407074_407074 ; 
   reg __407074_407074;
   reg _407075_407075 ; 
   reg __407075_407075;
   reg _407076_407076 ; 
   reg __407076_407076;
   reg _407077_407077 ; 
   reg __407077_407077;
   reg _407078_407078 ; 
   reg __407078_407078;
   reg _407079_407079 ; 
   reg __407079_407079;
   reg _407080_407080 ; 
   reg __407080_407080;
   reg _407081_407081 ; 
   reg __407081_407081;
   reg _407082_407082 ; 
   reg __407082_407082;
   reg _407083_407083 ; 
   reg __407083_407083;
   reg _407084_407084 ; 
   reg __407084_407084;
   reg _407085_407085 ; 
   reg __407085_407085;
   reg _407086_407086 ; 
   reg __407086_407086;
   reg _407087_407087 ; 
   reg __407087_407087;
   reg _407088_407088 ; 
   reg __407088_407088;
   reg _407089_407089 ; 
   reg __407089_407089;
   reg _407090_407090 ; 
   reg __407090_407090;
   reg _407091_407091 ; 
   reg __407091_407091;
   reg _407092_407092 ; 
   reg __407092_407092;
   reg _407093_407093 ; 
   reg __407093_407093;
   reg _407094_407094 ; 
   reg __407094_407094;
   reg _407095_407095 ; 
   reg __407095_407095;
   reg _407096_407096 ; 
   reg __407096_407096;
   reg _407097_407097 ; 
   reg __407097_407097;
   reg _407098_407098 ; 
   reg __407098_407098;
   reg _407099_407099 ; 
   reg __407099_407099;
   reg _407100_407100 ; 
   reg __407100_407100;
   reg _407101_407101 ; 
   reg __407101_407101;
   reg _407102_407102 ; 
   reg __407102_407102;
   reg _407103_407103 ; 
   reg __407103_407103;
   reg _407104_407104 ; 
   reg __407104_407104;
   reg _407105_407105 ; 
   reg __407105_407105;
   reg _407106_407106 ; 
   reg __407106_407106;
   reg _407107_407107 ; 
   reg __407107_407107;
   reg _407108_407108 ; 
   reg __407108_407108;
   reg _407109_407109 ; 
   reg __407109_407109;
   reg _407110_407110 ; 
   reg __407110_407110;
   reg _407111_407111 ; 
   reg __407111_407111;
   reg _407112_407112 ; 
   reg __407112_407112;
   reg _407113_407113 ; 
   reg __407113_407113;
   reg _407114_407114 ; 
   reg __407114_407114;
   reg _407115_407115 ; 
   reg __407115_407115;
   reg _407116_407116 ; 
   reg __407116_407116;
   reg _407117_407117 ; 
   reg __407117_407117;
   reg _407118_407118 ; 
   reg __407118_407118;
   reg _407119_407119 ; 
   reg __407119_407119;
   reg _407120_407120 ; 
   reg __407120_407120;
   reg _407121_407121 ; 
   reg __407121_407121;
   reg _407122_407122 ; 
   reg __407122_407122;
   reg _407123_407123 ; 
   reg __407123_407123;
   reg _407124_407124 ; 
   reg __407124_407124;
   reg _407125_407125 ; 
   reg __407125_407125;
   reg _407126_407126 ; 
   reg __407126_407126;
   reg _407127_407127 ; 
   reg __407127_407127;
   reg _407128_407128 ; 
   reg __407128_407128;
   reg _407129_407129 ; 
   reg __407129_407129;
   reg _407130_407130 ; 
   reg __407130_407130;
   reg _407131_407131 ; 
   reg __407131_407131;
   reg _407132_407132 ; 
   reg __407132_407132;
   reg _407133_407133 ; 
   reg __407133_407133;
   reg _407134_407134 ; 
   reg __407134_407134;
   reg _407135_407135 ; 
   reg __407135_407135;
   reg _407136_407136 ; 
   reg __407136_407136;
   reg _407137_407137 ; 
   reg __407137_407137;
   reg _407138_407138 ; 
   reg __407138_407138;
   reg _407139_407139 ; 
   reg __407139_407139;
   reg _407140_407140 ; 
   reg __407140_407140;
   reg _407141_407141 ; 
   reg __407141_407141;
   reg _407142_407142 ; 
   reg __407142_407142;
   reg _407143_407143 ; 
   reg __407143_407143;
   reg _407144_407144 ; 
   reg __407144_407144;
   reg _407145_407145 ; 
   reg __407145_407145;
   reg _407146_407146 ; 
   reg __407146_407146;
   reg _407147_407147 ; 
   reg __407147_407147;
   reg _407148_407148 ; 
   reg __407148_407148;
   reg _407149_407149 ; 
   reg __407149_407149;
   reg _407150_407150 ; 
   reg __407150_407150;
   reg _407151_407151 ; 
   reg __407151_407151;
   reg _407152_407152 ; 
   reg __407152_407152;
   reg _407153_407153 ; 
   reg __407153_407153;
   reg _407154_407154 ; 
   reg __407154_407154;
   reg _407155_407155 ; 
   reg __407155_407155;
   reg _407156_407156 ; 
   reg __407156_407156;
   reg _407157_407157 ; 
   reg __407157_407157;
   reg _407158_407158 ; 
   reg __407158_407158;
   reg _407159_407159 ; 
   reg __407159_407159;
   reg _407160_407160 ; 
   reg __407160_407160;
   reg _407161_407161 ; 
   reg __407161_407161;
   reg _407162_407162 ; 
   reg __407162_407162;
   reg _407163_407163 ; 
   reg __407163_407163;
   reg _407164_407164 ; 
   reg __407164_407164;
   reg _407165_407165 ; 
   reg __407165_407165;
   reg _407166_407166 ; 
   reg __407166_407166;
   reg _407167_407167 ; 
   reg __407167_407167;
   reg _407168_407168 ; 
   reg __407168_407168;
   reg _407169_407169 ; 
   reg __407169_407169;
   reg _407170_407170 ; 
   reg __407170_407170;
   reg _407171_407171 ; 
   reg __407171_407171;
   reg _407172_407172 ; 
   reg __407172_407172;
   reg _407173_407173 ; 
   reg __407173_407173;
   reg _407174_407174 ; 
   reg __407174_407174;
   reg _407175_407175 ; 
   reg __407175_407175;
   reg _407176_407176 ; 
   reg __407176_407176;
   reg _407177_407177 ; 
   reg __407177_407177;
   reg _407178_407178 ; 
   reg __407178_407178;
   reg _407179_407179 ; 
   reg __407179_407179;
   reg _407180_407180 ; 
   reg __407180_407180;
   reg _407181_407181 ; 
   reg __407181_407181;
   reg _407182_407182 ; 
   reg __407182_407182;
   reg _407183_407183 ; 
   reg __407183_407183;
   reg _407184_407184 ; 
   reg __407184_407184;
   reg _407185_407185 ; 
   reg __407185_407185;
   reg _407186_407186 ; 
   reg __407186_407186;
   reg _407187_407187 ; 
   reg __407187_407187;
   reg _407188_407188 ; 
   reg __407188_407188;
   reg _407189_407189 ; 
   reg __407189_407189;
   reg _407190_407190 ; 
   reg __407190_407190;
   reg _407191_407191 ; 
   reg __407191_407191;
   reg _407192_407192 ; 
   reg __407192_407192;
   reg _407193_407193 ; 
   reg __407193_407193;
   reg _407194_407194 ; 
   reg __407194_407194;
   reg _407195_407195 ; 
   reg __407195_407195;
   reg _407196_407196 ; 
   reg __407196_407196;
   reg _407197_407197 ; 
   reg __407197_407197;
   reg _407198_407198 ; 
   reg __407198_407198;
   reg _407199_407199 ; 
   reg __407199_407199;
   reg _407200_407200 ; 
   reg __407200_407200;
   reg _407201_407201 ; 
   reg __407201_407201;
   reg _407202_407202 ; 
   reg __407202_407202;
   reg _407203_407203 ; 
   reg __407203_407203;
   reg _407204_407204 ; 
   reg __407204_407204;
   reg _407205_407205 ; 
   reg __407205_407205;
   reg _407206_407206 ; 
   reg __407206_407206;
   reg _407207_407207 ; 
   reg __407207_407207;
   reg _407208_407208 ; 
   reg __407208_407208;
   reg _407209_407209 ; 
   reg __407209_407209;
   reg _407210_407210 ; 
   reg __407210_407210;
   reg _407211_407211 ; 
   reg __407211_407211;
   reg _407212_407212 ; 
   reg __407212_407212;
   reg _407213_407213 ; 
   reg __407213_407213;
   reg _407214_407214 ; 
   reg __407214_407214;
   reg _407215_407215 ; 
   reg __407215_407215;
   reg _407216_407216 ; 
   reg __407216_407216;
   reg _407217_407217 ; 
   reg __407217_407217;
   reg _407218_407218 ; 
   reg __407218_407218;
   reg _407219_407219 ; 
   reg __407219_407219;
   reg _407220_407220 ; 
   reg __407220_407220;
   reg _407221_407221 ; 
   reg __407221_407221;
   reg _407222_407222 ; 
   reg __407222_407222;
   reg _407223_407223 ; 
   reg __407223_407223;
   reg _407224_407224 ; 
   reg __407224_407224;
   reg _407225_407225 ; 
   reg __407225_407225;
   reg _407226_407226 ; 
   reg __407226_407226;
   reg _407227_407227 ; 
   reg __407227_407227;
   reg _407228_407228 ; 
   reg __407228_407228;
   reg _407229_407229 ; 
   reg __407229_407229;
   reg _407230_407230 ; 
   reg __407230_407230;
   reg _407231_407231 ; 
   reg __407231_407231;
   reg _407232_407232 ; 
   reg __407232_407232;
   reg _407233_407233 ; 
   reg __407233_407233;
   reg _407234_407234 ; 
   reg __407234_407234;
   reg _407235_407235 ; 
   reg __407235_407235;
   reg _407236_407236 ; 
   reg __407236_407236;
   reg _407237_407237 ; 
   reg __407237_407237;
   reg _407238_407238 ; 
   reg __407238_407238;
   reg _407239_407239 ; 
   reg __407239_407239;
   reg _407240_407240 ; 
   reg __407240_407240;
   reg _407241_407241 ; 
   reg __407241_407241;
   reg _407242_407242 ; 
   reg __407242_407242;
   reg _407243_407243 ; 
   reg __407243_407243;
   reg _407244_407244 ; 
   reg __407244_407244;
   reg _407245_407245 ; 
   reg __407245_407245;
   reg _407246_407246 ; 
   reg __407246_407246;
   reg _407247_407247 ; 
   reg __407247_407247;
   reg _407248_407248 ; 
   reg __407248_407248;
   reg _407249_407249 ; 
   reg __407249_407249;
   reg _407250_407250 ; 
   reg __407250_407250;
   reg _407251_407251 ; 
   reg __407251_407251;
   reg _407252_407252 ; 
   reg __407252_407252;
   reg _407253_407253 ; 
   reg __407253_407253;
   reg _407254_407254 ; 
   reg __407254_407254;
   reg _407255_407255 ; 
   reg __407255_407255;
   reg _407256_407256 ; 
   reg __407256_407256;
   reg _407257_407257 ; 
   reg __407257_407257;
   reg _407258_407258 ; 
   reg __407258_407258;
   reg _407259_407259 ; 
   reg __407259_407259;
   reg _407260_407260 ; 
   reg __407260_407260;
   reg _407261_407261 ; 
   reg __407261_407261;
   reg _407262_407262 ; 
   reg __407262_407262;
   reg _407263_407263 ; 
   reg __407263_407263;
   reg _407264_407264 ; 
   reg __407264_407264;
   reg _407265_407265 ; 
   reg __407265_407265;
   reg _407266_407266 ; 
   reg __407266_407266;
   reg _407267_407267 ; 
   reg __407267_407267;
   reg _407268_407268 ; 
   reg __407268_407268;
   reg _407269_407269 ; 
   reg __407269_407269;
   reg _407270_407270 ; 
   reg __407270_407270;
   reg _407271_407271 ; 
   reg __407271_407271;
   reg _407272_407272 ; 
   reg __407272_407272;
   reg _407273_407273 ; 
   reg __407273_407273;
   reg _407274_407274 ; 
   reg __407274_407274;
   reg _407275_407275 ; 
   reg __407275_407275;
   reg _407276_407276 ; 
   reg __407276_407276;
   reg _407277_407277 ; 
   reg __407277_407277;
   reg _407278_407278 ; 
   reg __407278_407278;
   reg _407279_407279 ; 
   reg __407279_407279;
   reg _407280_407280 ; 
   reg __407280_407280;
   reg _407281_407281 ; 
   reg __407281_407281;
   reg _407282_407282 ; 
   reg __407282_407282;
   reg _407283_407283 ; 
   reg __407283_407283;
   reg _407284_407284 ; 
   reg __407284_407284;
   reg _407285_407285 ; 
   reg __407285_407285;
   reg _407286_407286 ; 
   reg __407286_407286;
   reg _407287_407287 ; 
   reg __407287_407287;
   reg _407288_407288 ; 
   reg __407288_407288;
   reg _407289_407289 ; 
   reg __407289_407289;
   reg _407290_407290 ; 
   reg __407290_407290;
   reg _407291_407291 ; 
   reg __407291_407291;
   reg _407292_407292 ; 
   reg __407292_407292;
   reg _407293_407293 ; 
   reg __407293_407293;
   reg _407294_407294 ; 
   reg __407294_407294;
   reg _407295_407295 ; 
   reg __407295_407295;
   reg _407296_407296 ; 
   reg __407296_407296;
   reg _407297_407297 ; 
   reg __407297_407297;
   reg _407298_407298 ; 
   reg __407298_407298;
   reg _407299_407299 ; 
   reg __407299_407299;
   reg _407300_407300 ; 
   reg __407300_407300;
   reg _407301_407301 ; 
   reg __407301_407301;
   reg _407302_407302 ; 
   reg __407302_407302;
   reg _407303_407303 ; 
   reg __407303_407303;
   reg _407304_407304 ; 
   reg __407304_407304;
   reg _407305_407305 ; 
   reg __407305_407305;
   reg _407306_407306 ; 
   reg __407306_407306;
   reg _407307_407307 ; 
   reg __407307_407307;
   reg _407308_407308 ; 
   reg __407308_407308;
   reg _407309_407309 ; 
   reg __407309_407309;
   reg _407310_407310 ; 
   reg __407310_407310;
   reg _407311_407311 ; 
   reg __407311_407311;
   reg _407312_407312 ; 
   reg __407312_407312;
   reg _407313_407313 ; 
   reg __407313_407313;
   reg _407314_407314 ; 
   reg __407314_407314;
   reg _407315_407315 ; 
   reg __407315_407315;
   reg _407316_407316 ; 
   reg __407316_407316;
   reg _407317_407317 ; 
   reg __407317_407317;
   reg _407318_407318 ; 
   reg __407318_407318;
   reg _407319_407319 ; 
   reg __407319_407319;
   reg _407320_407320 ; 
   reg __407320_407320;
   reg _407321_407321 ; 
   reg __407321_407321;
   reg _407322_407322 ; 
   reg __407322_407322;
   reg _407323_407323 ; 
   reg __407323_407323;
   reg _407324_407324 ; 
   reg __407324_407324;
   reg _407325_407325 ; 
   reg __407325_407325;
   reg _407326_407326 ; 
   reg __407326_407326;
   reg _407327_407327 ; 
   reg __407327_407327;
   reg _407328_407328 ; 
   reg __407328_407328;
   reg _407329_407329 ; 
   reg __407329_407329;
   reg _407330_407330 ; 
   reg __407330_407330;
   reg _407331_407331 ; 
   reg __407331_407331;
   reg _407332_407332 ; 
   reg __407332_407332;
   reg _407333_407333 ; 
   reg __407333_407333;
   reg _407334_407334 ; 
   reg __407334_407334;
   reg _407335_407335 ; 
   reg __407335_407335;
   reg _407336_407336 ; 
   reg __407336_407336;
   reg _407337_407337 ; 
   reg __407337_407337;
   reg _407338_407338 ; 
   reg __407338_407338;
   reg _407339_407339 ; 
   reg __407339_407339;
   reg _407340_407340 ; 
   reg __407340_407340;
   reg _407341_407341 ; 
   reg __407341_407341;
   reg _407342_407342 ; 
   reg __407342_407342;
   reg _407343_407343 ; 
   reg __407343_407343;
   reg _407344_407344 ; 
   reg __407344_407344;
   reg _407345_407345 ; 
   reg __407345_407345;
   reg _407346_407346 ; 
   reg __407346_407346;
   reg _407347_407347 ; 
   reg __407347_407347;
   reg _407348_407348 ; 
   reg __407348_407348;
   reg _407349_407349 ; 
   reg __407349_407349;
   reg _407350_407350 ; 
   reg __407350_407350;
   reg _407351_407351 ; 
   reg __407351_407351;
   reg _407352_407352 ; 
   reg __407352_407352;
   reg _407353_407353 ; 
   reg __407353_407353;
   reg _407354_407354 ; 
   reg __407354_407354;
   reg _407355_407355 ; 
   reg __407355_407355;
   reg _407356_407356 ; 
   reg __407356_407356;
   reg _407357_407357 ; 
   reg __407357_407357;
   reg _407358_407358 ; 
   reg __407358_407358;
   reg _407359_407359 ; 
   reg __407359_407359;
   reg _407360_407360 ; 
   reg __407360_407360;
   reg _407361_407361 ; 
   reg __407361_407361;
   reg _407362_407362 ; 
   reg __407362_407362;
   reg _407363_407363 ; 
   reg __407363_407363;
   reg _407364_407364 ; 
   reg __407364_407364;
   reg _407365_407365 ; 
   reg __407365_407365;
   reg _407366_407366 ; 
   reg __407366_407366;
   reg _407367_407367 ; 
   reg __407367_407367;
   reg _407368_407368 ; 
   reg __407368_407368;
   reg _407369_407369 ; 
   reg __407369_407369;
   reg _407370_407370 ; 
   reg __407370_407370;
   reg _407371_407371 ; 
   reg __407371_407371;
   reg _407372_407372 ; 
   reg __407372_407372;
   reg _407373_407373 ; 
   reg __407373_407373;
   reg _407374_407374 ; 
   reg __407374_407374;
   reg _407375_407375 ; 
   reg __407375_407375;
   reg _407376_407376 ; 
   reg __407376_407376;
   reg _407377_407377 ; 
   reg __407377_407377;
   reg _407378_407378 ; 
   reg __407378_407378;
   reg _407379_407379 ; 
   reg __407379_407379;
   reg _407380_407380 ; 
   reg __407380_407380;
   reg _407381_407381 ; 
   reg __407381_407381;
   reg _407382_407382 ; 
   reg __407382_407382;
   reg _407383_407383 ; 
   reg __407383_407383;
   reg _407384_407384 ; 
   reg __407384_407384;
   reg _407385_407385 ; 
   reg __407385_407385;
   reg _407386_407386 ; 
   reg __407386_407386;
   reg _407387_407387 ; 
   reg __407387_407387;
   reg _407388_407388 ; 
   reg __407388_407388;
   reg _407389_407389 ; 
   reg __407389_407389;
   reg _407390_407390 ; 
   reg __407390_407390;
   reg _407391_407391 ; 
   reg __407391_407391;
   reg _407392_407392 ; 
   reg __407392_407392;
   reg _407393_407393 ; 
   reg __407393_407393;
   reg _407394_407394 ; 
   reg __407394_407394;
   reg _407395_407395 ; 
   reg __407395_407395;
   reg _407396_407396 ; 
   reg __407396_407396;
   reg _407397_407397 ; 
   reg __407397_407397;
   reg _407398_407398 ; 
   reg __407398_407398;
   reg _407399_407399 ; 
   reg __407399_407399;
   reg _407400_407400 ; 
   reg __407400_407400;
   reg _407401_407401 ; 
   reg __407401_407401;
   reg _407402_407402 ; 
   reg __407402_407402;
   reg _407403_407403 ; 
   reg __407403_407403;
   reg _407404_407404 ; 
   reg __407404_407404;
   reg _407405_407405 ; 
   reg __407405_407405;
   reg _407406_407406 ; 
   reg __407406_407406;
   reg _407407_407407 ; 
   reg __407407_407407;
   reg _407408_407408 ; 
   reg __407408_407408;
   reg _407409_407409 ; 
   reg __407409_407409;
   reg _407410_407410 ; 
   reg __407410_407410;
   reg _407411_407411 ; 
   reg __407411_407411;
   reg _407412_407412 ; 
   reg __407412_407412;
   reg _407413_407413 ; 
   reg __407413_407413;
   reg _407414_407414 ; 
   reg __407414_407414;
   reg _407415_407415 ; 
   reg __407415_407415;
   reg _407416_407416 ; 
   reg __407416_407416;
   reg _407417_407417 ; 
   reg __407417_407417;
   reg _407418_407418 ; 
   reg __407418_407418;
   reg _407419_407419 ; 
   reg __407419_407419;
   reg _407420_407420 ; 
   reg __407420_407420;
   reg _407421_407421 ; 
   reg __407421_407421;
   reg _407422_407422 ; 
   reg __407422_407422;
   reg _407423_407423 ; 
   reg __407423_407423;
   reg _407424_407424 ; 
   reg __407424_407424;
   reg _407425_407425 ; 
   reg __407425_407425;
   reg _407426_407426 ; 
   reg __407426_407426;
   reg _407427_407427 ; 
   reg __407427_407427;
   reg _407428_407428 ; 
   reg __407428_407428;
   reg _407429_407429 ; 
   reg __407429_407429;
   reg _407430_407430 ; 
   reg __407430_407430;
   reg _407431_407431 ; 
   reg __407431_407431;
   reg _407432_407432 ; 
   reg __407432_407432;
   reg _407433_407433 ; 
   reg __407433_407433;
   reg _407434_407434 ; 
   reg __407434_407434;
   reg _407435_407435 ; 
   reg __407435_407435;
   reg _407436_407436 ; 
   reg __407436_407436;
   reg _407437_407437 ; 
   reg __407437_407437;
   reg _407438_407438 ; 
   reg __407438_407438;
   reg _407439_407439 ; 
   reg __407439_407439;
   reg _407440_407440 ; 
   reg __407440_407440;
   reg _407441_407441 ; 
   reg __407441_407441;
   reg _407442_407442 ; 
   reg __407442_407442;
   reg _407443_407443 ; 
   reg __407443_407443;
   reg _407444_407444 ; 
   reg __407444_407444;
   reg _407445_407445 ; 
   reg __407445_407445;
   reg _407446_407446 ; 
   reg __407446_407446;
   reg _407447_407447 ; 
   reg __407447_407447;
   reg _407448_407448 ; 
   reg __407448_407448;
   reg _407449_407449 ; 
   reg __407449_407449;
   reg _407450_407450 ; 
   reg __407450_407450;
   reg _407451_407451 ; 
   reg __407451_407451;
   reg _407452_407452 ; 
   reg __407452_407452;
   reg _407453_407453 ; 
   reg __407453_407453;
   reg _407454_407454 ; 
   reg __407454_407454;
   reg _407455_407455 ; 
   reg __407455_407455;
   reg _407456_407456 ; 
   reg __407456_407456;
   reg _407457_407457 ; 
   reg __407457_407457;
   reg _407458_407458 ; 
   reg __407458_407458;
   reg _407459_407459 ; 
   reg __407459_407459;
   reg _407460_407460 ; 
   reg __407460_407460;
   reg _407461_407461 ; 
   reg __407461_407461;
   reg _407462_407462 ; 
   reg __407462_407462;
   reg _407463_407463 ; 
   reg __407463_407463;
   reg _407464_407464 ; 
   reg __407464_407464;
   reg _407465_407465 ; 
   reg __407465_407465;
   reg _407466_407466 ; 
   reg __407466_407466;
   reg _407467_407467 ; 
   reg __407467_407467;
   reg _407468_407468 ; 
   reg __407468_407468;
   reg _407469_407469 ; 
   reg __407469_407469;
   reg _407470_407470 ; 
   reg __407470_407470;
   reg _407471_407471 ; 
   reg __407471_407471;
   reg _407472_407472 ; 
   reg __407472_407472;
   reg _407473_407473 ; 
   reg __407473_407473;
   reg _407474_407474 ; 
   reg __407474_407474;
   reg _407475_407475 ; 
   reg __407475_407475;
   reg _407476_407476 ; 
   reg __407476_407476;
   reg _407477_407477 ; 
   reg __407477_407477;
   reg _407478_407478 ; 
   reg __407478_407478;
   reg _407479_407479 ; 
   reg __407479_407479;
   reg _407480_407480 ; 
   reg __407480_407480;
   reg _407481_407481 ; 
   reg __407481_407481;
   reg _407482_407482 ; 
   reg __407482_407482;
   reg _407483_407483 ; 
   reg __407483_407483;
   reg _407484_407484 ; 
   reg __407484_407484;
   reg _407485_407485 ; 
   reg __407485_407485;
   reg _407486_407486 ; 
   reg __407486_407486;
   reg _407487_407487 ; 
   reg __407487_407487;
   reg _407488_407488 ; 
   reg __407488_407488;
   reg _407489_407489 ; 
   reg __407489_407489;
   reg _407490_407490 ; 
   reg __407490_407490;
   reg _407491_407491 ; 
   reg __407491_407491;
   reg _407492_407492 ; 
   reg __407492_407492;
   reg _407493_407493 ; 
   reg __407493_407493;
   reg _407494_407494 ; 
   reg __407494_407494;
   reg _407495_407495 ; 
   reg __407495_407495;
   reg _407496_407496 ; 
   reg __407496_407496;
   reg _407497_407497 ; 
   reg __407497_407497;
   reg _407498_407498 ; 
   reg __407498_407498;
   reg _407499_407499 ; 
   reg __407499_407499;
   reg _407500_407500 ; 
   reg __407500_407500;
   reg _407501_407501 ; 
   reg __407501_407501;
   reg _407502_407502 ; 
   reg __407502_407502;
   reg _407503_407503 ; 
   reg __407503_407503;
   reg _407504_407504 ; 
   reg __407504_407504;
   reg _407505_407505 ; 
   reg __407505_407505;
   reg _407506_407506 ; 
   reg __407506_407506;
   reg _407507_407507 ; 
   reg __407507_407507;
   reg _407508_407508 ; 
   reg __407508_407508;
   reg _407509_407509 ; 
   reg __407509_407509;
   reg _407510_407510 ; 
   reg __407510_407510;
   reg _407511_407511 ; 
   reg __407511_407511;
   reg _407512_407512 ; 
   reg __407512_407512;
   reg _407513_407513 ; 
   reg __407513_407513;
   reg _407514_407514 ; 
   reg __407514_407514;
   reg _407515_407515 ; 
   reg __407515_407515;
   reg _407516_407516 ; 
   reg __407516_407516;
   reg _407517_407517 ; 
   reg __407517_407517;
   reg _407518_407518 ; 
   reg __407518_407518;
   reg _407519_407519 ; 
   reg __407519_407519;
   reg _407520_407520 ; 
   reg __407520_407520;
   reg _407521_407521 ; 
   reg __407521_407521;
   reg _407522_407522 ; 
   reg __407522_407522;
   reg _407523_407523 ; 
   reg __407523_407523;
   reg _407524_407524 ; 
   reg __407524_407524;
   reg _407525_407525 ; 
   reg __407525_407525;
   reg _407526_407526 ; 
   reg __407526_407526;
   reg _407527_407527 ; 
   reg __407527_407527;
   reg _407528_407528 ; 
   reg __407528_407528;
   reg _407529_407529 ; 
   reg __407529_407529;
   reg _407530_407530 ; 
   reg __407530_407530;
   reg _407531_407531 ; 
   reg __407531_407531;
   reg _407532_407532 ; 
   reg __407532_407532;
   reg _407533_407533 ; 
   reg __407533_407533;
   reg _407534_407534 ; 
   reg __407534_407534;
   reg _407535_407535 ; 
   reg __407535_407535;
   reg _407536_407536 ; 
   reg __407536_407536;
   reg _407537_407537 ; 
   reg __407537_407537;
   reg _407538_407538 ; 
   reg __407538_407538;
   reg _407539_407539 ; 
   reg __407539_407539;
   reg _407540_407540 ; 
   reg __407540_407540;
   reg _407541_407541 ; 
   reg __407541_407541;
   reg _407542_407542 ; 
   reg __407542_407542;
   reg _407543_407543 ; 
   reg __407543_407543;
   reg _407544_407544 ; 
   reg __407544_407544;
   reg _407545_407545 ; 
   reg __407545_407545;
   reg _407546_407546 ; 
   reg __407546_407546;
   reg _407547_407547 ; 
   reg __407547_407547;
   reg _407548_407548 ; 
   reg __407548_407548;
   reg _407549_407549 ; 
   reg __407549_407549;
   reg _407550_407550 ; 
   reg __407550_407550;
   reg _407551_407551 ; 
   reg __407551_407551;
   reg _407552_407552 ; 
   reg __407552_407552;
   reg _407553_407553 ; 
   reg __407553_407553;
   reg _407554_407554 ; 
   reg __407554_407554;
   reg _407555_407555 ; 
   reg __407555_407555;
   reg _407556_407556 ; 
   reg __407556_407556;
   reg _407557_407557 ; 
   reg __407557_407557;
   reg _407558_407558 ; 
   reg __407558_407558;
   reg _407559_407559 ; 
   reg __407559_407559;
   reg _407560_407560 ; 
   reg __407560_407560;
   reg _407561_407561 ; 
   reg __407561_407561;
   reg _407562_407562 ; 
   reg __407562_407562;
   reg _407563_407563 ; 
   reg __407563_407563;
   reg _407564_407564 ; 
   reg __407564_407564;
   reg _407565_407565 ; 
   reg __407565_407565;
   reg _407566_407566 ; 
   reg __407566_407566;
   reg _407567_407567 ; 
   reg __407567_407567;
   reg _407568_407568 ; 
   reg __407568_407568;
   reg _407569_407569 ; 
   reg __407569_407569;
   reg _407570_407570 ; 
   reg __407570_407570;
   reg _407571_407571 ; 
   reg __407571_407571;
   reg _407572_407572 ; 
   reg __407572_407572;
   reg _407573_407573 ; 
   reg __407573_407573;
   reg _407574_407574 ; 
   reg __407574_407574;
   reg _407575_407575 ; 
   reg __407575_407575;
   reg _407576_407576 ; 
   reg __407576_407576;
   reg _407577_407577 ; 
   reg __407577_407577;
   reg _407578_407578 ; 
   reg __407578_407578;
   reg _407579_407579 ; 
   reg __407579_407579;
   reg _407580_407580 ; 
   reg __407580_407580;
   reg _407581_407581 ; 
   reg __407581_407581;
   reg _407582_407582 ; 
   reg __407582_407582;
   reg _407583_407583 ; 
   reg __407583_407583;
   reg _407584_407584 ; 
   reg __407584_407584;
   reg _407585_407585 ; 
   reg __407585_407585;
   reg _407586_407586 ; 
   reg __407586_407586;
   reg _407587_407587 ; 
   reg __407587_407587;
   reg _407588_407588 ; 
   reg __407588_407588;
   reg _407589_407589 ; 
   reg __407589_407589;
   reg _407590_407590 ; 
   reg __407590_407590;
   reg _407591_407591 ; 
   reg __407591_407591;
   reg _407592_407592 ; 
   reg __407592_407592;
   reg _407593_407593 ; 
   reg __407593_407593;
   reg _407594_407594 ; 
   reg __407594_407594;
   reg _407595_407595 ; 
   reg __407595_407595;
   reg _407596_407596 ; 
   reg __407596_407596;
   reg _407597_407597 ; 
   reg __407597_407597;
   reg _407598_407598 ; 
   reg __407598_407598;
   reg _407599_407599 ; 
   reg __407599_407599;
   reg _407600_407600 ; 
   reg __407600_407600;
   reg _407601_407601 ; 
   reg __407601_407601;
   reg _407602_407602 ; 
   reg __407602_407602;
   reg _407603_407603 ; 
   reg __407603_407603;
   reg _407604_407604 ; 
   reg __407604_407604;
   reg _407605_407605 ; 
   reg __407605_407605;
   reg _407606_407606 ; 
   reg __407606_407606;
   reg _407607_407607 ; 
   reg __407607_407607;
   reg _407608_407608 ; 
   reg __407608_407608;
   reg _407609_407609 ; 
   reg __407609_407609;
   reg _407610_407610 ; 
   reg __407610_407610;
   reg _407611_407611 ; 
   reg __407611_407611;
   reg _407612_407612 ; 
   reg __407612_407612;
   reg _407613_407613 ; 
   reg __407613_407613;
   reg _407614_407614 ; 
   reg __407614_407614;
   reg _407615_407615 ; 
   reg __407615_407615;
   reg _407616_407616 ; 
   reg __407616_407616;
   reg _407617_407617 ; 
   reg __407617_407617;
   reg _407618_407618 ; 
   reg __407618_407618;
   reg _407619_407619 ; 
   reg __407619_407619;
   reg _407620_407620 ; 
   reg __407620_407620;
   reg _407621_407621 ; 
   reg __407621_407621;
   reg _407622_407622 ; 
   reg __407622_407622;
   reg _407623_407623 ; 
   reg __407623_407623;
   reg _407624_407624 ; 
   reg __407624_407624;
   reg _407625_407625 ; 
   reg __407625_407625;
   reg _407626_407626 ; 
   reg __407626_407626;
   reg _407627_407627 ; 
   reg __407627_407627;
   reg _407628_407628 ; 
   reg __407628_407628;
   reg _407629_407629 ; 
   reg __407629_407629;
   reg _407630_407630 ; 
   reg __407630_407630;
   reg _407631_407631 ; 
   reg __407631_407631;
   reg _407632_407632 ; 
   reg __407632_407632;
   reg _407633_407633 ; 
   reg __407633_407633;
   reg _407634_407634 ; 
   reg __407634_407634;
   reg _407635_407635 ; 
   reg __407635_407635;
   reg _407636_407636 ; 
   reg __407636_407636;
   reg _407637_407637 ; 
   reg __407637_407637;
   reg _407638_407638 ; 
   reg __407638_407638;
   reg _407639_407639 ; 
   reg __407639_407639;
   reg _407640_407640 ; 
   reg __407640_407640;
   reg _407641_407641 ; 
   reg __407641_407641;
   reg _407642_407642 ; 
   reg __407642_407642;
   reg _407643_407643 ; 
   reg __407643_407643;
   reg _407644_407644 ; 
   reg __407644_407644;
   reg _407645_407645 ; 
   reg __407645_407645;
   reg _407646_407646 ; 
   reg __407646_407646;
   reg _407647_407647 ; 
   reg __407647_407647;
   reg _407648_407648 ; 
   reg __407648_407648;
   reg _407649_407649 ; 
   reg __407649_407649;
   reg _407650_407650 ; 
   reg __407650_407650;
   reg _407651_407651 ; 
   reg __407651_407651;
   reg _407652_407652 ; 
   reg __407652_407652;
   reg _407653_407653 ; 
   reg __407653_407653;
   reg _407654_407654 ; 
   reg __407654_407654;
   reg _407655_407655 ; 
   reg __407655_407655;
   reg _407656_407656 ; 
   reg __407656_407656;
   reg _407657_407657 ; 
   reg __407657_407657;
   reg _407658_407658 ; 
   reg __407658_407658;
   reg _407659_407659 ; 
   reg __407659_407659;
   reg _407660_407660 ; 
   reg __407660_407660;
   reg _407661_407661 ; 
   reg __407661_407661;
   reg _407662_407662 ; 
   reg __407662_407662;
   reg _407663_407663 ; 
   reg __407663_407663;
   reg _407664_407664 ; 
   reg __407664_407664;
   reg _407665_407665 ; 
   reg __407665_407665;
   reg _407666_407666 ; 
   reg __407666_407666;
   reg _407667_407667 ; 
   reg __407667_407667;
   reg _407668_407668 ; 
   reg __407668_407668;
   reg _407669_407669 ; 
   reg __407669_407669;
   reg _407670_407670 ; 
   reg __407670_407670;
   reg _407671_407671 ; 
   reg __407671_407671;
   reg _407672_407672 ; 
   reg __407672_407672;
   reg _407673_407673 ; 
   reg __407673_407673;
   reg _407674_407674 ; 
   reg __407674_407674;
   reg _407675_407675 ; 
   reg __407675_407675;
   reg _407676_407676 ; 
   reg __407676_407676;
   reg _407677_407677 ; 
   reg __407677_407677;
   reg _407678_407678 ; 
   reg __407678_407678;
   reg _407679_407679 ; 
   reg __407679_407679;
   reg _407680_407680 ; 
   reg __407680_407680;
   reg _407681_407681 ; 
   reg __407681_407681;
   reg _407682_407682 ; 
   reg __407682_407682;
   reg _407683_407683 ; 
   reg __407683_407683;
   reg _407684_407684 ; 
   reg __407684_407684;
   reg _407685_407685 ; 
   reg __407685_407685;
   reg _407686_407686 ; 
   reg __407686_407686;
   reg _407687_407687 ; 
   reg __407687_407687;
   reg _407688_407688 ; 
   reg __407688_407688;
   reg _407689_407689 ; 
   reg __407689_407689;
   reg _407690_407690 ; 
   reg __407690_407690;
   reg _407691_407691 ; 
   reg __407691_407691;
   reg _407692_407692 ; 
   reg __407692_407692;
   reg _407693_407693 ; 
   reg __407693_407693;
   reg _407694_407694 ; 
   reg __407694_407694;
   reg _407695_407695 ; 
   reg __407695_407695;
   reg _407696_407696 ; 
   reg __407696_407696;
   reg _407697_407697 ; 
   reg __407697_407697;
   reg _407698_407698 ; 
   reg __407698_407698;
   reg _407699_407699 ; 
   reg __407699_407699;
   reg _407700_407700 ; 
   reg __407700_407700;
   reg _407701_407701 ; 
   reg __407701_407701;
   reg _407702_407702 ; 
   reg __407702_407702;
   reg _407703_407703 ; 
   reg __407703_407703;
   reg _407704_407704 ; 
   reg __407704_407704;
   reg _407705_407705 ; 
   reg __407705_407705;
   reg _407706_407706 ; 
   reg __407706_407706;
   reg _407707_407707 ; 
   reg __407707_407707;
   reg _407708_407708 ; 
   reg __407708_407708;
   reg _407709_407709 ; 
   reg __407709_407709;
   reg _407710_407710 ; 
   reg __407710_407710;
   reg _407711_407711 ; 
   reg __407711_407711;
   reg _407712_407712 ; 
   reg __407712_407712;
   reg _407713_407713 ; 
   reg __407713_407713;
   reg _407714_407714 ; 
   reg __407714_407714;
   reg _407715_407715 ; 
   reg __407715_407715;
   reg _407716_407716 ; 
   reg __407716_407716;
   reg _407717_407717 ; 
   reg __407717_407717;
   reg _407718_407718 ; 
   reg __407718_407718;
   reg _407719_407719 ; 
   reg __407719_407719;
   reg _407720_407720 ; 
   reg __407720_407720;
   reg _407721_407721 ; 
   reg __407721_407721;
   reg _407722_407722 ; 
   reg __407722_407722;
   reg _407723_407723 ; 
   reg __407723_407723;
   reg _407724_407724 ; 
   reg __407724_407724;
   reg _407725_407725 ; 
   reg __407725_407725;
   reg _407726_407726 ; 
   reg __407726_407726;
   reg _407727_407727 ; 
   reg __407727_407727;
   reg _407728_407728 ; 
   reg __407728_407728;
   reg _407729_407729 ; 
   reg __407729_407729;
   reg _407730_407730 ; 
   reg __407730_407730;
   reg _407731_407731 ; 
   reg __407731_407731;
   reg _407732_407732 ; 
   reg __407732_407732;
   reg _407733_407733 ; 
   reg __407733_407733;
   reg _407734_407734 ; 
   reg __407734_407734;
   reg _407735_407735 ; 
   reg __407735_407735;
   reg _407736_407736 ; 
   reg __407736_407736;
   reg _407737_407737 ; 
   reg __407737_407737;
   reg _407738_407738 ; 
   reg __407738_407738;
   reg _407739_407739 ; 
   reg __407739_407739;
   reg _407740_407740 ; 
   reg __407740_407740;
   reg _407741_407741 ; 
   reg __407741_407741;
   reg _407742_407742 ; 
   reg __407742_407742;
   reg _407743_407743 ; 
   reg __407743_407743;
   reg _407744_407744 ; 
   reg __407744_407744;
   reg _407745_407745 ; 
   reg __407745_407745;
   reg _407746_407746 ; 
   reg __407746_407746;
   reg _407747_407747 ; 
   reg __407747_407747;
   reg _407748_407748 ; 
   reg __407748_407748;
   reg _407749_407749 ; 
   reg __407749_407749;
   reg _407750_407750 ; 
   reg __407750_407750;
   reg _407751_407751 ; 
   reg __407751_407751;
   reg _407752_407752 ; 
   reg __407752_407752;
   reg _407753_407753 ; 
   reg __407753_407753;
   reg _407754_407754 ; 
   reg __407754_407754;
   reg _407755_407755 ; 
   reg __407755_407755;
   reg _407756_407756 ; 
   reg __407756_407756;
   reg _407757_407757 ; 
   reg __407757_407757;
   reg _407758_407758 ; 
   reg __407758_407758;
   reg _407759_407759 ; 
   reg __407759_407759;
   reg _407760_407760 ; 
   reg __407760_407760;
   reg _407761_407761 ; 
   reg __407761_407761;
   reg _407762_407762 ; 
   reg __407762_407762;
   reg _407763_407763 ; 
   reg __407763_407763;
   reg _407764_407764 ; 
   reg __407764_407764;
   reg _407765_407765 ; 
   reg __407765_407765;
   reg _407766_407766 ; 
   reg __407766_407766;
   reg _407767_407767 ; 
   reg __407767_407767;
   reg _407768_407768 ; 
   reg __407768_407768;
   reg _407769_407769 ; 
   reg __407769_407769;
   reg _407770_407770 ; 
   reg __407770_407770;
   reg _407771_407771 ; 
   reg __407771_407771;
   reg _407772_407772 ; 
   reg __407772_407772;
   reg _407773_407773 ; 
   reg __407773_407773;
   reg _407774_407774 ; 
   reg __407774_407774;
   reg _407775_407775 ; 
   reg __407775_407775;
   reg _407776_407776 ; 
   reg __407776_407776;
   reg _407777_407777 ; 
   reg __407777_407777;
   reg _407778_407778 ; 
   reg __407778_407778;
   reg _407779_407779 ; 
   reg __407779_407779;
   reg _407780_407780 ; 
   reg __407780_407780;
   reg _407781_407781 ; 
   reg __407781_407781;
   reg _407782_407782 ; 
   reg __407782_407782;
   reg _407783_407783 ; 
   reg __407783_407783;
   reg _407784_407784 ; 
   reg __407784_407784;
   reg _407785_407785 ; 
   reg __407785_407785;
   reg _407786_407786 ; 
   reg __407786_407786;
   reg _407787_407787 ; 
   reg __407787_407787;
   reg _407788_407788 ; 
   reg __407788_407788;
   reg _407789_407789 ; 
   reg __407789_407789;
   reg _407790_407790 ; 
   reg __407790_407790;
   reg _407791_407791 ; 
   reg __407791_407791;
   reg _407792_407792 ; 
   reg __407792_407792;
   reg _407793_407793 ; 
   reg __407793_407793;
   reg _407794_407794 ; 
   reg __407794_407794;
   reg _407795_407795 ; 
   reg __407795_407795;
   reg _407796_407796 ; 
   reg __407796_407796;
   reg _407797_407797 ; 
   reg __407797_407797;
   reg _407798_407798 ; 
   reg __407798_407798;
   reg _407799_407799 ; 
   reg __407799_407799;
   reg _407800_407800 ; 
   reg __407800_407800;
   reg _407801_407801 ; 
   reg __407801_407801;
   reg _407802_407802 ; 
   reg __407802_407802;
   reg _407803_407803 ; 
   reg __407803_407803;
   reg _407804_407804 ; 
   reg __407804_407804;
   reg _407805_407805 ; 
   reg __407805_407805;
   reg _407806_407806 ; 
   reg __407806_407806;
   reg _407807_407807 ; 
   reg __407807_407807;
   reg _407808_407808 ; 
   reg __407808_407808;
   reg _407809_407809 ; 
   reg __407809_407809;
   reg _407810_407810 ; 
   reg __407810_407810;
   reg _407811_407811 ; 
   reg __407811_407811;
   reg _407812_407812 ; 
   reg __407812_407812;
   reg _407813_407813 ; 
   reg __407813_407813;
   reg _407814_407814 ; 
   reg __407814_407814;
   reg _407815_407815 ; 
   reg __407815_407815;
   reg _407816_407816 ; 
   reg __407816_407816;
   reg _407817_407817 ; 
   reg __407817_407817;
   reg _407818_407818 ; 
   reg __407818_407818;
   reg _407819_407819 ; 
   reg __407819_407819;
   reg _407820_407820 ; 
   reg __407820_407820;
   reg _407821_407821 ; 
   reg __407821_407821;
   reg _407822_407822 ; 
   reg __407822_407822;
   reg _407823_407823 ; 
   reg __407823_407823;
   reg _407824_407824 ; 
   reg __407824_407824;
   reg _407825_407825 ; 
   reg __407825_407825;
   reg _407826_407826 ; 
   reg __407826_407826;
   reg _407827_407827 ; 
   reg __407827_407827;
   reg _407828_407828 ; 
   reg __407828_407828;
   reg _407829_407829 ; 
   reg __407829_407829;
   reg _407830_407830 ; 
   reg __407830_407830;
   reg _407831_407831 ; 
   reg __407831_407831;
   reg _407832_407832 ; 
   reg __407832_407832;
   reg _407833_407833 ; 
   reg __407833_407833;
   reg _407834_407834 ; 
   reg __407834_407834;
   reg _407835_407835 ; 
   reg __407835_407835;
   reg _407836_407836 ; 
   reg __407836_407836;
   reg _407837_407837 ; 
   reg __407837_407837;
   reg _407838_407838 ; 
   reg __407838_407838;
   reg _407839_407839 ; 
   reg __407839_407839;
   reg _407840_407840 ; 
   reg __407840_407840;
   reg _407841_407841 ; 
   reg __407841_407841;
   reg _407842_407842 ; 
   reg __407842_407842;
   reg _407843_407843 ; 
   reg __407843_407843;
   reg _407844_407844 ; 
   reg __407844_407844;
   reg _407845_407845 ; 
   reg __407845_407845;
   reg _407846_407846 ; 
   reg __407846_407846;
   reg _407847_407847 ; 
   reg __407847_407847;
   reg _407848_407848 ; 
   reg __407848_407848;
   reg _407849_407849 ; 
   reg __407849_407849;
   reg _407850_407850 ; 
   reg __407850_407850;
   reg _407851_407851 ; 
   reg __407851_407851;
   reg _407852_407852 ; 
   reg __407852_407852;
   reg _407853_407853 ; 
   reg __407853_407853;
   reg _407854_407854 ; 
   reg __407854_407854;
   reg _407855_407855 ; 
   reg __407855_407855;
   reg _407856_407856 ; 
   reg __407856_407856;
   reg _407857_407857 ; 
   reg __407857_407857;
   reg _407858_407858 ; 
   reg __407858_407858;
   reg _407859_407859 ; 
   reg __407859_407859;
   reg _407860_407860 ; 
   reg __407860_407860;
   reg _407861_407861 ; 
   reg __407861_407861;
   reg _407862_407862 ; 
   reg __407862_407862;
   reg _407863_407863 ; 
   reg __407863_407863;
   reg _407864_407864 ; 
   reg __407864_407864;
   reg _407865_407865 ; 
   reg __407865_407865;
   reg _407866_407866 ; 
   reg __407866_407866;
   reg _407867_407867 ; 
   reg __407867_407867;
   reg _407868_407868 ; 
   reg __407868_407868;
   reg _407869_407869 ; 
   reg __407869_407869;
   reg _407870_407870 ; 
   reg __407870_407870;
   reg _407871_407871 ; 
   reg __407871_407871;
   reg _407872_407872 ; 
   reg __407872_407872;
   reg _407873_407873 ; 
   reg __407873_407873;
   reg _407874_407874 ; 
   reg __407874_407874;
   reg _407875_407875 ; 
   reg __407875_407875;
   reg _407876_407876 ; 
   reg __407876_407876;
   reg _407877_407877 ; 
   reg __407877_407877;
   reg _407878_407878 ; 
   reg __407878_407878;
   reg _407879_407879 ; 
   reg __407879_407879;
   reg _407880_407880 ; 
   reg __407880_407880;
   reg _407881_407881 ; 
   reg __407881_407881;
   reg _407882_407882 ; 
   reg __407882_407882;
   reg _407883_407883 ; 
   reg __407883_407883;
   reg _407884_407884 ; 
   reg __407884_407884;
   reg _407885_407885 ; 
   reg __407885_407885;
   reg _407886_407886 ; 
   reg __407886_407886;
   reg _407887_407887 ; 
   reg __407887_407887;
   reg _407888_407888 ; 
   reg __407888_407888;
   reg _407889_407889 ; 
   reg __407889_407889;
   reg _407890_407890 ; 
   reg __407890_407890;
   reg _407891_407891 ; 
   reg __407891_407891;
   reg _407892_407892 ; 
   reg __407892_407892;
   reg _407893_407893 ; 
   reg __407893_407893;
   reg _407894_407894 ; 
   reg __407894_407894;
   reg _407895_407895 ; 
   reg __407895_407895;
   reg _407896_407896 ; 
   reg __407896_407896;
   reg _407897_407897 ; 
   reg __407897_407897;
   reg _407898_407898 ; 
   reg __407898_407898;
   reg _407899_407899 ; 
   reg __407899_407899;
   reg _407900_407900 ; 
   reg __407900_407900;
   reg _407901_407901 ; 
   reg __407901_407901;
   reg _407902_407902 ; 
   reg __407902_407902;
   reg _407903_407903 ; 
   reg __407903_407903;
   reg _407904_407904 ; 
   reg __407904_407904;
   reg _407905_407905 ; 
   reg __407905_407905;
   reg _407906_407906 ; 
   reg __407906_407906;
   reg _407907_407907 ; 
   reg __407907_407907;
   reg _407908_407908 ; 
   reg __407908_407908;
   reg _407909_407909 ; 
   reg __407909_407909;
   reg _407910_407910 ; 
   reg __407910_407910;
   reg _407911_407911 ; 
   reg __407911_407911;
   reg _407912_407912 ; 
   reg __407912_407912;
   reg _407913_407913 ; 
   reg __407913_407913;
   reg _407914_407914 ; 
   reg __407914_407914;
   reg _407915_407915 ; 
   reg __407915_407915;
   reg _407916_407916 ; 
   reg __407916_407916;
   reg _407917_407917 ; 
   reg __407917_407917;
   reg _407918_407918 ; 
   reg __407918_407918;
   reg _407919_407919 ; 
   reg __407919_407919;
   reg _407920_407920 ; 
   reg __407920_407920;
   reg _407921_407921 ; 
   reg __407921_407921;
   reg _407922_407922 ; 
   reg __407922_407922;
   reg _407923_407923 ; 
   reg __407923_407923;
   reg _407924_407924 ; 
   reg __407924_407924;
   reg _407925_407925 ; 
   reg __407925_407925;
   reg _407926_407926 ; 
   reg __407926_407926;
   reg _407927_407927 ; 
   reg __407927_407927;
   reg _407928_407928 ; 
   reg __407928_407928;
   reg _407929_407929 ; 
   reg __407929_407929;
   reg _407930_407930 ; 
   reg __407930_407930;
   reg _407931_407931 ; 
   reg __407931_407931;
   reg _407932_407932 ; 
   reg __407932_407932;
   reg _407933_407933 ; 
   reg __407933_407933;
   reg _407934_407934 ; 
   reg __407934_407934;
   reg _407935_407935 ; 
   reg __407935_407935;
   reg _407936_407936 ; 
   reg __407936_407936;
   reg _407937_407937 ; 
   reg __407937_407937;
   reg _407938_407938 ; 
   reg __407938_407938;
   reg _407939_407939 ; 
   reg __407939_407939;
   reg _407940_407940 ; 
   reg __407940_407940;
   reg _407941_407941 ; 
   reg __407941_407941;
   reg _407942_407942 ; 
   reg __407942_407942;
   reg _407943_407943 ; 
   reg __407943_407943;
   reg _407944_407944 ; 
   reg __407944_407944;
   reg _407945_407945 ; 
   reg __407945_407945;
   reg _407946_407946 ; 
   reg __407946_407946;
   reg _407947_407947 ; 
   reg __407947_407947;
   reg _407948_407948 ; 
   reg __407948_407948;
   reg _407949_407949 ; 
   reg __407949_407949;
   reg _407950_407950 ; 
   reg __407950_407950;
   reg _407951_407951 ; 
   reg __407951_407951;
   reg _407952_407952 ; 
   reg __407952_407952;
   reg _407953_407953 ; 
   reg __407953_407953;
   reg _407954_407954 ; 
   reg __407954_407954;
   reg _407955_407955 ; 
   reg __407955_407955;
   reg _407956_407956 ; 
   reg __407956_407956;
   reg _407957_407957 ; 
   reg __407957_407957;
   reg _407958_407958 ; 
   reg __407958_407958;
   reg _407959_407959 ; 
   reg __407959_407959;
   reg _407960_407960 ; 
   reg __407960_407960;
   reg _407961_407961 ; 
   reg __407961_407961;
   reg _407962_407962 ; 
   reg __407962_407962;
   reg _407963_407963 ; 
   reg __407963_407963;
   reg _407964_407964 ; 
   reg __407964_407964;
   reg _407965_407965 ; 
   reg __407965_407965;
   reg _407966_407966 ; 
   reg __407966_407966;
   reg _407967_407967 ; 
   reg __407967_407967;
   reg _407968_407968 ; 
   reg __407968_407968;
   reg _407969_407969 ; 
   reg __407969_407969;
   reg _407970_407970 ; 
   reg __407970_407970;
   reg _407971_407971 ; 
   reg __407971_407971;
   reg _407972_407972 ; 
   reg __407972_407972;
   reg _407973_407973 ; 
   reg __407973_407973;
   reg _407974_407974 ; 
   reg __407974_407974;
   reg _407975_407975 ; 
   reg __407975_407975;
   reg _407976_407976 ; 
   reg __407976_407976;
   reg _407977_407977 ; 
   reg __407977_407977;
   reg _407978_407978 ; 
   reg __407978_407978;
   reg _407979_407979 ; 
   reg __407979_407979;
   reg _407980_407980 ; 
   reg __407980_407980;
   reg _407981_407981 ; 
   reg __407981_407981;
   reg _407982_407982 ; 
   reg __407982_407982;
   reg _407983_407983 ; 
   reg __407983_407983;
   reg _407984_407984 ; 
   reg __407984_407984;
   reg _407985_407985 ; 
   reg __407985_407985;
   reg _407986_407986 ; 
   reg __407986_407986;
   reg _407987_407987 ; 
   reg __407987_407987;
   reg _407988_407988 ; 
   reg __407988_407988;
   reg _407989_407989 ; 
   reg __407989_407989;
   reg _407990_407990 ; 
   reg __407990_407990;
   reg _407991_407991 ; 
   reg __407991_407991;
   reg _407992_407992 ; 
   reg __407992_407992;
   reg _407993_407993 ; 
   reg __407993_407993;
   reg _407994_407994 ; 
   reg __407994_407994;
   reg _407995_407995 ; 
   reg __407995_407995;
   reg _407996_407996 ; 
   reg __407996_407996;
   reg _407997_407997 ; 
   reg __407997_407997;
   reg _407998_407998 ; 
   reg __407998_407998;
   reg _407999_407999 ; 
   reg __407999_407999;
   reg _408000_408000 ; 
   reg __408000_408000;
   reg _408001_408001 ; 
   reg __408001_408001;
   reg _408002_408002 ; 
   reg __408002_408002;
   reg _408003_408003 ; 
   reg __408003_408003;
   reg _408004_408004 ; 
   reg __408004_408004;
   reg _408005_408005 ; 
   reg __408005_408005;
   reg _408006_408006 ; 
   reg __408006_408006;
   reg _408007_408007 ; 
   reg __408007_408007;
   reg _408008_408008 ; 
   reg __408008_408008;
   reg _408009_408009 ; 
   reg __408009_408009;
   reg _408010_408010 ; 
   reg __408010_408010;
   reg _408011_408011 ; 
   reg __408011_408011;
   reg _408012_408012 ; 
   reg __408012_408012;
   reg _408013_408013 ; 
   reg __408013_408013;
   reg _408014_408014 ; 
   reg __408014_408014;
   reg _408015_408015 ; 
   reg __408015_408015;
   reg _408016_408016 ; 
   reg __408016_408016;
   reg _408017_408017 ; 
   reg __408017_408017;
   reg _408018_408018 ; 
   reg __408018_408018;
   reg _408019_408019 ; 
   reg __408019_408019;
   reg _408020_408020 ; 
   reg __408020_408020;
   reg _408021_408021 ; 
   reg __408021_408021;
   reg _408022_408022 ; 
   reg __408022_408022;
   reg _408023_408023 ; 
   reg __408023_408023;
   reg _408024_408024 ; 
   reg __408024_408024;
   reg _408025_408025 ; 
   reg __408025_408025;
   reg _408026_408026 ; 
   reg __408026_408026;
   reg _408027_408027 ; 
   reg __408027_408027;
   reg _408028_408028 ; 
   reg __408028_408028;
   reg _408029_408029 ; 
   reg __408029_408029;
   reg _408030_408030 ; 
   reg __408030_408030;
   reg _408031_408031 ; 
   reg __408031_408031;
   reg _408032_408032 ; 
   reg __408032_408032;
   reg _408033_408033 ; 
   reg __408033_408033;
   reg _408034_408034 ; 
   reg __408034_408034;
   reg _408035_408035 ; 
   reg __408035_408035;
   reg _408036_408036 ; 
   reg __408036_408036;
   reg _408037_408037 ; 
   reg __408037_408037;
   reg _408038_408038 ; 
   reg __408038_408038;
   reg _408039_408039 ; 
   reg __408039_408039;
   reg _408040_408040 ; 
   reg __408040_408040;
   reg _408041_408041 ; 
   reg __408041_408041;
   reg _408042_408042 ; 
   reg __408042_408042;
   reg _408043_408043 ; 
   reg __408043_408043;
   reg _408044_408044 ; 
   reg __408044_408044;
   reg _408045_408045 ; 
   reg __408045_408045;
   reg _408046_408046 ; 
   reg __408046_408046;
   reg _408047_408047 ; 
   reg __408047_408047;
   reg _408048_408048 ; 
   reg __408048_408048;
   reg _408049_408049 ; 
   reg __408049_408049;
   reg _408050_408050 ; 
   reg __408050_408050;
   reg _408051_408051 ; 
   reg __408051_408051;
   reg _408052_408052 ; 
   reg __408052_408052;
   reg _408053_408053 ; 
   reg __408053_408053;
   reg _408054_408054 ; 
   reg __408054_408054;
   reg _408055_408055 ; 
   reg __408055_408055;
   reg _408056_408056 ; 
   reg __408056_408056;
   reg _408057_408057 ; 
   reg __408057_408057;
   reg _408058_408058 ; 
   reg __408058_408058;
   reg _408059_408059 ; 
   reg __408059_408059;
   reg _408060_408060 ; 
   reg __408060_408060;
   reg _408061_408061 ; 
   reg __408061_408061;
   reg _408062_408062 ; 
   reg __408062_408062;
   reg _408063_408063 ; 
   reg __408063_408063;
   reg _408064_408064 ; 
   reg __408064_408064;
   reg _408065_408065 ; 
   reg __408065_408065;
   reg _408066_408066 ; 
   reg __408066_408066;
   reg _408067_408067 ; 
   reg __408067_408067;
   reg _408068_408068 ; 
   reg __408068_408068;
   reg _408069_408069 ; 
   reg __408069_408069;
   reg _408070_408070 ; 
   reg __408070_408070;
   reg _408071_408071 ; 
   reg __408071_408071;
   reg _408072_408072 ; 
   reg __408072_408072;
   reg _408073_408073 ; 
   reg __408073_408073;
   reg _408074_408074 ; 
   reg __408074_408074;
   reg _408075_408075 ; 
   reg __408075_408075;
   reg _408076_408076 ; 
   reg __408076_408076;
   reg _408077_408077 ; 
   reg __408077_408077;
   reg _408078_408078 ; 
   reg __408078_408078;
   reg _408079_408079 ; 
   reg __408079_408079;
   reg _408080_408080 ; 
   reg __408080_408080;
   reg _408081_408081 ; 
   reg __408081_408081;
   reg _408082_408082 ; 
   reg __408082_408082;
   reg _408083_408083 ; 
   reg __408083_408083;
   reg _408084_408084 ; 
   reg __408084_408084;
   reg _408085_408085 ; 
   reg __408085_408085;
   reg _408086_408086 ; 
   reg __408086_408086;
   reg _408087_408087 ; 
   reg __408087_408087;
   reg _408088_408088 ; 
   reg __408088_408088;
   reg _408089_408089 ; 
   reg __408089_408089;
   reg _408090_408090 ; 
   reg __408090_408090;
   reg _408091_408091 ; 
   reg __408091_408091;
   reg _408092_408092 ; 
   reg __408092_408092;
   reg _408093_408093 ; 
   reg __408093_408093;
   reg _408094_408094 ; 
   reg __408094_408094;
   reg _408095_408095 ; 
   reg __408095_408095;
   reg _408096_408096 ; 
   reg __408096_408096;
   reg _408097_408097 ; 
   reg __408097_408097;
   reg _408098_408098 ; 
   reg __408098_408098;
   reg _408099_408099 ; 
   reg __408099_408099;
   reg _408100_408100 ; 
   reg __408100_408100;
   reg _408101_408101 ; 
   reg __408101_408101;
   reg _408102_408102 ; 
   reg __408102_408102;
   reg _408103_408103 ; 
   reg __408103_408103;
   reg _408104_408104 ; 
   reg __408104_408104;
   reg _408105_408105 ; 
   reg __408105_408105;
   reg _408106_408106 ; 
   reg __408106_408106;
   reg _408107_408107 ; 
   reg __408107_408107;
   reg _408108_408108 ; 
   reg __408108_408108;
   reg _408109_408109 ; 
   reg __408109_408109;
   reg _408110_408110 ; 
   reg __408110_408110;
   reg _408111_408111 ; 
   reg __408111_408111;
   reg _408112_408112 ; 
   reg __408112_408112;
   reg _408113_408113 ; 
   reg __408113_408113;
   reg _408114_408114 ; 
   reg __408114_408114;
   reg _408115_408115 ; 
   reg __408115_408115;
   reg _408116_408116 ; 
   reg __408116_408116;
   reg _408117_408117 ; 
   reg __408117_408117;
   reg _408118_408118 ; 
   reg __408118_408118;
   reg _408119_408119 ; 
   reg __408119_408119;
   reg _408120_408120 ; 
   reg __408120_408120;
   reg _408121_408121 ; 
   reg __408121_408121;
   reg _408122_408122 ; 
   reg __408122_408122;
   reg _408123_408123 ; 
   reg __408123_408123;
   reg _408124_408124 ; 
   reg __408124_408124;
   reg _408125_408125 ; 
   reg __408125_408125;
   reg _408126_408126 ; 
   reg __408126_408126;
   reg _408127_408127 ; 
   reg __408127_408127;
   reg _408128_408128 ; 
   reg __408128_408128;
   reg _408129_408129 ; 
   reg __408129_408129;
   reg _408130_408130 ; 
   reg __408130_408130;
   reg _408131_408131 ; 
   reg __408131_408131;
   reg _408132_408132 ; 
   reg __408132_408132;
   reg _408133_408133 ; 
   reg __408133_408133;
   reg _408134_408134 ; 
   reg __408134_408134;
   reg _408135_408135 ; 
   reg __408135_408135;
   reg _408136_408136 ; 
   reg __408136_408136;
   reg _408137_408137 ; 
   reg __408137_408137;
   reg _408138_408138 ; 
   reg __408138_408138;
   reg _408139_408139 ; 
   reg __408139_408139;
   reg _408140_408140 ; 
   reg __408140_408140;
   reg _408141_408141 ; 
   reg __408141_408141;
   reg _408142_408142 ; 
   reg __408142_408142;
   reg _408143_408143 ; 
   reg __408143_408143;
   reg _408144_408144 ; 
   reg __408144_408144;
   reg _408145_408145 ; 
   reg __408145_408145;
   reg _408146_408146 ; 
   reg __408146_408146;
   reg _408147_408147 ; 
   reg __408147_408147;
   reg _408148_408148 ; 
   reg __408148_408148;
   reg _408149_408149 ; 
   reg __408149_408149;
   reg _408150_408150 ; 
   reg __408150_408150;
   reg _408151_408151 ; 
   reg __408151_408151;
   reg _408152_408152 ; 
   reg __408152_408152;
   reg _408153_408153 ; 
   reg __408153_408153;
   reg _408154_408154 ; 
   reg __408154_408154;
   reg _408155_408155 ; 
   reg __408155_408155;
   reg _408156_408156 ; 
   reg __408156_408156;
   reg _408157_408157 ; 
   reg __408157_408157;
   reg _408158_408158 ; 
   reg __408158_408158;
   reg _408159_408159 ; 
   reg __408159_408159;
   reg _408160_408160 ; 
   reg __408160_408160;
   reg _408161_408161 ; 
   reg __408161_408161;
   reg _408162_408162 ; 
   reg __408162_408162;
   reg _408163_408163 ; 
   reg __408163_408163;
   reg _408164_408164 ; 
   reg __408164_408164;
   reg _408165_408165 ; 
   reg __408165_408165;
   reg _408166_408166 ; 
   reg __408166_408166;
   reg _408167_408167 ; 
   reg __408167_408167;
   reg _408168_408168 ; 
   reg __408168_408168;
   reg _408169_408169 ; 
   reg __408169_408169;
   reg _408170_408170 ; 
   reg __408170_408170;
   reg _408171_408171 ; 
   reg __408171_408171;
   reg _408172_408172 ; 
   reg __408172_408172;
   reg _408173_408173 ; 
   reg __408173_408173;
   reg _408174_408174 ; 
   reg __408174_408174;
   reg _408175_408175 ; 
   reg __408175_408175;
   reg _408176_408176 ; 
   reg __408176_408176;
   reg _408177_408177 ; 
   reg __408177_408177;
   reg _408178_408178 ; 
   reg __408178_408178;
   reg _408179_408179 ; 
   reg __408179_408179;
   reg _408180_408180 ; 
   reg __408180_408180;
   reg _408181_408181 ; 
   reg __408181_408181;
   reg _408182_408182 ; 
   reg __408182_408182;
   reg _408183_408183 ; 
   reg __408183_408183;
   reg _408184_408184 ; 
   reg __408184_408184;
   reg _408185_408185 ; 
   reg __408185_408185;
   reg _408186_408186 ; 
   reg __408186_408186;
   reg _408187_408187 ; 
   reg __408187_408187;
   reg _408188_408188 ; 
   reg __408188_408188;
   reg _408189_408189 ; 
   reg __408189_408189;
   reg _408190_408190 ; 
   reg __408190_408190;
   reg _408191_408191 ; 
   reg __408191_408191;
   reg _408192_408192 ; 
   reg __408192_408192;
   reg _408193_408193 ; 
   reg __408193_408193;
   reg _408194_408194 ; 
   reg __408194_408194;
   reg _408195_408195 ; 
   reg __408195_408195;
   reg _408196_408196 ; 
   reg __408196_408196;
   reg _408197_408197 ; 
   reg __408197_408197;
   reg _408198_408198 ; 
   reg __408198_408198;
   reg _408199_408199 ; 
   reg __408199_408199;
   reg _408200_408200 ; 
   reg __408200_408200;
   reg _408201_408201 ; 
   reg __408201_408201;
   reg _408202_408202 ; 
   reg __408202_408202;
   reg _408203_408203 ; 
   reg __408203_408203;
   reg _408204_408204 ; 
   reg __408204_408204;
   reg _408205_408205 ; 
   reg __408205_408205;
   reg _408206_408206 ; 
   reg __408206_408206;
   reg _408207_408207 ; 
   reg __408207_408207;
   reg _408208_408208 ; 
   reg __408208_408208;
   reg _408209_408209 ; 
   reg __408209_408209;
   reg _408210_408210 ; 
   reg __408210_408210;
   reg _408211_408211 ; 
   reg __408211_408211;
   reg _408212_408212 ; 
   reg __408212_408212;
   reg _408213_408213 ; 
   reg __408213_408213;
   reg _408214_408214 ; 
   reg __408214_408214;
   reg _408215_408215 ; 
   reg __408215_408215;
   reg _408216_408216 ; 
   reg __408216_408216;
   reg _408217_408217 ; 
   reg __408217_408217;
   reg _408218_408218 ; 
   reg __408218_408218;
   reg _408219_408219 ; 
   reg __408219_408219;
   reg _408220_408220 ; 
   reg __408220_408220;
   reg _408221_408221 ; 
   reg __408221_408221;
   reg _408222_408222 ; 
   reg __408222_408222;
   reg _408223_408223 ; 
   reg __408223_408223;
   reg _408224_408224 ; 
   reg __408224_408224;
   reg _408225_408225 ; 
   reg __408225_408225;
   reg _408226_408226 ; 
   reg __408226_408226;
   reg _408227_408227 ; 
   reg __408227_408227;
   reg _408228_408228 ; 
   reg __408228_408228;
   reg _408229_408229 ; 
   reg __408229_408229;
   reg _408230_408230 ; 
   reg __408230_408230;
   reg _408231_408231 ; 
   reg __408231_408231;
   reg _408232_408232 ; 
   reg __408232_408232;
   reg _408233_408233 ; 
   reg __408233_408233;
   reg _408234_408234 ; 
   reg __408234_408234;
   reg _408235_408235 ; 
   reg __408235_408235;
   reg _408236_408236 ; 
   reg __408236_408236;
   reg _408237_408237 ; 
   reg __408237_408237;
   reg _408238_408238 ; 
   reg __408238_408238;
   reg _408239_408239 ; 
   reg __408239_408239;
   reg _408240_408240 ; 
   reg __408240_408240;
   reg _408241_408241 ; 
   reg __408241_408241;
   reg _408242_408242 ; 
   reg __408242_408242;
   reg _408243_408243 ; 
   reg __408243_408243;
   reg _408244_408244 ; 
   reg __408244_408244;
   reg _408245_408245 ; 
   reg __408245_408245;
   reg _408246_408246 ; 
   reg __408246_408246;
   reg _408247_408247 ; 
   reg __408247_408247;
   reg _408248_408248 ; 
   reg __408248_408248;
   reg _408249_408249 ; 
   reg __408249_408249;
   reg _408250_408250 ; 
   reg __408250_408250;
   reg _408251_408251 ; 
   reg __408251_408251;
   reg _408252_408252 ; 
   reg __408252_408252;
   reg _408253_408253 ; 
   reg __408253_408253;
   reg _408254_408254 ; 
   reg __408254_408254;
   reg _408255_408255 ; 
   reg __408255_408255;
   reg _408256_408256 ; 
   reg __408256_408256;
   reg _408257_408257 ; 
   reg __408257_408257;
   reg _408258_408258 ; 
   reg __408258_408258;
   reg _408259_408259 ; 
   reg __408259_408259;
   reg _408260_408260 ; 
   reg __408260_408260;
   reg _408261_408261 ; 
   reg __408261_408261;
   reg _408262_408262 ; 
   reg __408262_408262;
   reg _408263_408263 ; 
   reg __408263_408263;
   reg _408264_408264 ; 
   reg __408264_408264;
   reg _408265_408265 ; 
   reg __408265_408265;
   reg _408266_408266 ; 
   reg __408266_408266;
   reg _408267_408267 ; 
   reg __408267_408267;
   reg _408268_408268 ; 
   reg __408268_408268;
   reg _408269_408269 ; 
   reg __408269_408269;
   reg _408270_408270 ; 
   reg __408270_408270;
   reg _408271_408271 ; 
   reg __408271_408271;
   reg _408272_408272 ; 
   reg __408272_408272;
   reg _408273_408273 ; 
   reg __408273_408273;
   reg _408274_408274 ; 
   reg __408274_408274;
   reg _408275_408275 ; 
   reg __408275_408275;
   reg _408276_408276 ; 
   reg __408276_408276;
   reg _408277_408277 ; 
   reg __408277_408277;
   reg _408278_408278 ; 
   reg __408278_408278;
   reg _408279_408279 ; 
   reg __408279_408279;
   reg _408280_408280 ; 
   reg __408280_408280;
   reg _408281_408281 ; 
   reg __408281_408281;
   reg _408282_408282 ; 
   reg __408282_408282;
   reg _408283_408283 ; 
   reg __408283_408283;
   reg _408284_408284 ; 
   reg __408284_408284;
   reg _408285_408285 ; 
   reg __408285_408285;
   reg _408286_408286 ; 
   reg __408286_408286;
   reg _408287_408287 ; 
   reg __408287_408287;
   reg _408288_408288 ; 
   reg __408288_408288;
   reg _408289_408289 ; 
   reg __408289_408289;
   reg _408290_408290 ; 
   reg __408290_408290;
   reg _408291_408291 ; 
   reg __408291_408291;
   reg _408292_408292 ; 
   reg __408292_408292;
   reg _408293_408293 ; 
   reg __408293_408293;
   reg _408294_408294 ; 
   reg __408294_408294;
   reg _408295_408295 ; 
   reg __408295_408295;
   reg _408296_408296 ; 
   reg __408296_408296;
   reg _408297_408297 ; 
   reg __408297_408297;
   reg _408298_408298 ; 
   reg __408298_408298;
   reg _408299_408299 ; 
   reg __408299_408299;
   reg _408300_408300 ; 
   reg __408300_408300;
   reg _408301_408301 ; 
   reg __408301_408301;
   reg _408302_408302 ; 
   reg __408302_408302;
   reg _408303_408303 ; 
   reg __408303_408303;
   reg _408304_408304 ; 
   reg __408304_408304;
   reg _408305_408305 ; 
   reg __408305_408305;
   reg _408306_408306 ; 
   reg __408306_408306;
   reg _408307_408307 ; 
   reg __408307_408307;
   reg _408308_408308 ; 
   reg __408308_408308;
   reg _408309_408309 ; 
   reg __408309_408309;
   reg _408310_408310 ; 
   reg __408310_408310;
   reg _408311_408311 ; 
   reg __408311_408311;
   reg _408312_408312 ; 
   reg __408312_408312;
   reg _408313_408313 ; 
   reg __408313_408313;
   reg _408314_408314 ; 
   reg __408314_408314;
   reg _408315_408315 ; 
   reg __408315_408315;
   reg _408316_408316 ; 
   reg __408316_408316;
   reg _408317_408317 ; 
   reg __408317_408317;
   reg _408318_408318 ; 
   reg __408318_408318;
   reg _408319_408319 ; 
   reg __408319_408319;
   reg _408320_408320 ; 
   reg __408320_408320;
   reg _408321_408321 ; 
   reg __408321_408321;
   reg _408322_408322 ; 
   reg __408322_408322;
   reg _408323_408323 ; 
   reg __408323_408323;
   reg _408324_408324 ; 
   reg __408324_408324;
   reg _408325_408325 ; 
   reg __408325_408325;
   reg _408326_408326 ; 
   reg __408326_408326;
   reg _408327_408327 ; 
   reg __408327_408327;
   reg _408328_408328 ; 
   reg __408328_408328;
   reg _408329_408329 ; 
   reg __408329_408329;
   reg _408330_408330 ; 
   reg __408330_408330;
   reg _408331_408331 ; 
   reg __408331_408331;
   reg _408332_408332 ; 
   reg __408332_408332;
   reg _408333_408333 ; 
   reg __408333_408333;
   reg _408334_408334 ; 
   reg __408334_408334;
   reg _408335_408335 ; 
   reg __408335_408335;
   reg _408336_408336 ; 
   reg __408336_408336;
   reg _408337_408337 ; 
   reg __408337_408337;
   reg _408338_408338 ; 
   reg __408338_408338;
   reg _408339_408339 ; 
   reg __408339_408339;
   reg _408340_408340 ; 
   reg __408340_408340;
   reg _408341_408341 ; 
   reg __408341_408341;
   reg _408342_408342 ; 
   reg __408342_408342;
   reg _408343_408343 ; 
   reg __408343_408343;
   reg _408344_408344 ; 
   reg __408344_408344;
   reg _408345_408345 ; 
   reg __408345_408345;
   reg _408346_408346 ; 
   reg __408346_408346;
   reg _408347_408347 ; 
   reg __408347_408347;
   reg _408348_408348 ; 
   reg __408348_408348;
   reg _408349_408349 ; 
   reg __408349_408349;
   reg _408350_408350 ; 
   reg __408350_408350;
   reg _408351_408351 ; 
   reg __408351_408351;
   reg _408352_408352 ; 
   reg __408352_408352;
   reg _408353_408353 ; 
   reg __408353_408353;
   reg _408354_408354 ; 
   reg __408354_408354;
   reg _408355_408355 ; 
   reg __408355_408355;
   reg _408356_408356 ; 
   reg __408356_408356;
   reg _408357_408357 ; 
   reg __408357_408357;
   reg _408358_408358 ; 
   reg __408358_408358;
   reg _408359_408359 ; 
   reg __408359_408359;
   reg _408360_408360 ; 
   reg __408360_408360;
   reg _408361_408361 ; 
   reg __408361_408361;
   reg _408362_408362 ; 
   reg __408362_408362;
   reg _408363_408363 ; 
   reg __408363_408363;
   reg _408364_408364 ; 
   reg __408364_408364;
   reg _408365_408365 ; 
   reg __408365_408365;
   reg _408366_408366 ; 
   reg __408366_408366;
   reg _408367_408367 ; 
   reg __408367_408367;
   reg _408368_408368 ; 
   reg __408368_408368;
   reg _408369_408369 ; 
   reg __408369_408369;
   reg _408370_408370 ; 
   reg __408370_408370;
   reg _408371_408371 ; 
   reg __408371_408371;
   reg _408372_408372 ; 
   reg __408372_408372;
   reg _408373_408373 ; 
   reg __408373_408373;
   reg _408374_408374 ; 
   reg __408374_408374;
   reg _408375_408375 ; 
   reg __408375_408375;
   reg _408376_408376 ; 
   reg __408376_408376;
   reg _408377_408377 ; 
   reg __408377_408377;
   reg _408378_408378 ; 
   reg __408378_408378;
   reg _408379_408379 ; 
   reg __408379_408379;
   reg _408380_408380 ; 
   reg __408380_408380;
   reg _408381_408381 ; 
   reg __408381_408381;
   reg _408382_408382 ; 
   reg __408382_408382;
   reg _408383_408383 ; 
   reg __408383_408383;
   reg _408384_408384 ; 
   reg __408384_408384;
   reg _408385_408385 ; 
   reg __408385_408385;
   reg _408386_408386 ; 
   reg __408386_408386;
   reg _408387_408387 ; 
   reg __408387_408387;
   reg _408388_408388 ; 
   reg __408388_408388;
   reg _408389_408389 ; 
   reg __408389_408389;
   reg _408390_408390 ; 
   reg __408390_408390;
   reg _408391_408391 ; 
   reg __408391_408391;
   reg _408392_408392 ; 
   reg __408392_408392;
   reg _408393_408393 ; 
   reg __408393_408393;
   reg _408394_408394 ; 
   reg __408394_408394;
   reg _408395_408395 ; 
   reg __408395_408395;
   reg _408396_408396 ; 
   reg __408396_408396;
   reg _408397_408397 ; 
   reg __408397_408397;
   reg _408398_408398 ; 
   reg __408398_408398;
   reg _408399_408399 ; 
   reg __408399_408399;
   reg _408400_408400 ; 
   reg __408400_408400;
   reg _408401_408401 ; 
   reg __408401_408401;
   reg _408402_408402 ; 
   reg __408402_408402;
   reg _408403_408403 ; 
   reg __408403_408403;
   reg _408404_408404 ; 
   reg __408404_408404;
   reg _408405_408405 ; 
   reg __408405_408405;
   reg _408406_408406 ; 
   reg __408406_408406;
   reg _408407_408407 ; 
   reg __408407_408407;
   reg _408408_408408 ; 
   reg __408408_408408;
   reg _408409_408409 ; 
   reg __408409_408409;
   reg _408410_408410 ; 
   reg __408410_408410;
   reg _408411_408411 ; 
   reg __408411_408411;
   reg _408412_408412 ; 
   reg __408412_408412;
   reg _408413_408413 ; 
   reg __408413_408413;
   reg _408414_408414 ; 
   reg __408414_408414;
   reg _408415_408415 ; 
   reg __408415_408415;
   reg _408416_408416 ; 
   reg __408416_408416;
   reg _408417_408417 ; 
   reg __408417_408417;
   reg _408418_408418 ; 
   reg __408418_408418;
   reg _408419_408419 ; 
   reg __408419_408419;
   reg _408420_408420 ; 
   reg __408420_408420;
   reg _408421_408421 ; 
   reg __408421_408421;
   reg _408422_408422 ; 
   reg __408422_408422;
   reg _408423_408423 ; 
   reg __408423_408423;
   reg _408424_408424 ; 
   reg __408424_408424;
   reg _408425_408425 ; 
   reg __408425_408425;
   reg _408426_408426 ; 
   reg __408426_408426;
   reg _408427_408427 ; 
   reg __408427_408427;
   reg _408428_408428 ; 
   reg __408428_408428;
   reg _408429_408429 ; 
   reg __408429_408429;
   reg _408430_408430 ; 
   reg __408430_408430;
   reg _408431_408431 ; 
   reg __408431_408431;
   reg _408432_408432 ; 
   reg __408432_408432;
   reg _408433_408433 ; 
   reg __408433_408433;
   reg _408434_408434 ; 
   reg __408434_408434;
   reg _408435_408435 ; 
   reg __408435_408435;
   reg _408436_408436 ; 
   reg __408436_408436;
   reg _408437_408437 ; 
   reg __408437_408437;
   reg _408438_408438 ; 
   reg __408438_408438;
   reg _408439_408439 ; 
   reg __408439_408439;
   reg _408440_408440 ; 
   reg __408440_408440;
   reg _408441_408441 ; 
   reg __408441_408441;
   reg _408442_408442 ; 
   reg __408442_408442;
   reg _408443_408443 ; 
   reg __408443_408443;
   reg _408444_408444 ; 
   reg __408444_408444;
   reg _408445_408445 ; 
   reg __408445_408445;
   reg _408446_408446 ; 
   reg __408446_408446;
   reg _408447_408447 ; 
   reg __408447_408447;
   reg _408448_408448 ; 
   reg __408448_408448;
   reg _408449_408449 ; 
   reg __408449_408449;
   reg _408450_408450 ; 
   reg __408450_408450;
   reg _408451_408451 ; 
   reg __408451_408451;
   reg _408452_408452 ; 
   reg __408452_408452;
   reg _408453_408453 ; 
   reg __408453_408453;
   reg _408454_408454 ; 
   reg __408454_408454;
   reg _408455_408455 ; 
   reg __408455_408455;
   reg _408456_408456 ; 
   reg __408456_408456;
   reg _408457_408457 ; 
   reg __408457_408457;
   reg _408458_408458 ; 
   reg __408458_408458;
   reg _408459_408459 ; 
   reg __408459_408459;
   reg _408460_408460 ; 
   reg __408460_408460;
   reg _408461_408461 ; 
   reg __408461_408461;
   reg _408462_408462 ; 
   reg __408462_408462;
   reg _408463_408463 ; 
   reg __408463_408463;
   reg _408464_408464 ; 
   reg __408464_408464;
   reg _408465_408465 ; 
   reg __408465_408465;
   reg _408466_408466 ; 
   reg __408466_408466;
   reg _408467_408467 ; 
   reg __408467_408467;
   reg _408468_408468 ; 
   reg __408468_408468;
   reg _408469_408469 ; 
   reg __408469_408469;
   reg _408470_408470 ; 
   reg __408470_408470;
   reg _408471_408471 ; 
   reg __408471_408471;
   reg _408472_408472 ; 
   reg __408472_408472;
   reg _408473_408473 ; 
   reg __408473_408473;
   reg _408474_408474 ; 
   reg __408474_408474;
   reg _408475_408475 ; 
   reg __408475_408475;
   reg _408476_408476 ; 
   reg __408476_408476;
   reg _408477_408477 ; 
   reg __408477_408477;
   reg _408478_408478 ; 
   reg __408478_408478;
   reg _408479_408479 ; 
   reg __408479_408479;
   reg _408480_408480 ; 
   reg __408480_408480;
   reg _408481_408481 ; 
   reg __408481_408481;
   reg _408482_408482 ; 
   reg __408482_408482;
   reg _408483_408483 ; 
   reg __408483_408483;
   reg _408484_408484 ; 
   reg __408484_408484;
   reg _408485_408485 ; 
   reg __408485_408485;
   reg _408486_408486 ; 
   reg __408486_408486;
   reg _408487_408487 ; 
   reg __408487_408487;
   reg _408488_408488 ; 
   reg __408488_408488;
   reg _408489_408489 ; 
   reg __408489_408489;
   reg _408490_408490 ; 
   reg __408490_408490;
   reg _408491_408491 ; 
   reg __408491_408491;
   reg _408492_408492 ; 
   reg __408492_408492;
   reg _408493_408493 ; 
   reg __408493_408493;
   reg _408494_408494 ; 
   reg __408494_408494;
   reg _408495_408495 ; 
   reg __408495_408495;
   reg _408496_408496 ; 
   reg __408496_408496;
   reg _408497_408497 ; 
   reg __408497_408497;
   reg _408498_408498 ; 
   reg __408498_408498;
   reg _408499_408499 ; 
   reg __408499_408499;
   reg _408500_408500 ; 
   reg __408500_408500;
   reg _408501_408501 ; 
   reg __408501_408501;
   reg _408502_408502 ; 
   reg __408502_408502;
   reg _408503_408503 ; 
   reg __408503_408503;
   reg _408504_408504 ; 
   reg __408504_408504;
   reg _408505_408505 ; 
   reg __408505_408505;
   reg _408506_408506 ; 
   reg __408506_408506;
   reg _408507_408507 ; 
   reg __408507_408507;
   reg _408508_408508 ; 
   reg __408508_408508;
   reg _408509_408509 ; 
   reg __408509_408509;
   reg _408510_408510 ; 
   reg __408510_408510;
   reg _408511_408511 ; 
   reg __408511_408511;
   reg _408512_408512 ; 
   reg __408512_408512;
   reg _408513_408513 ; 
   reg __408513_408513;
   reg _408514_408514 ; 
   reg __408514_408514;
   reg _408515_408515 ; 
   reg __408515_408515;
   reg _408516_408516 ; 
   reg __408516_408516;
   reg _408517_408517 ; 
   reg __408517_408517;
   reg _408518_408518 ; 
   reg __408518_408518;
   reg _408519_408519 ; 
   reg __408519_408519;
   reg _408520_408520 ; 
   reg __408520_408520;
   reg _408521_408521 ; 
   reg __408521_408521;
   reg _408522_408522 ; 
   reg __408522_408522;
   reg _408523_408523 ; 
   reg __408523_408523;
   reg _408524_408524 ; 
   reg __408524_408524;
   reg _408525_408525 ; 
   reg __408525_408525;
   reg _408526_408526 ; 
   reg __408526_408526;
   reg _408527_408527 ; 
   reg __408527_408527;
   reg _408528_408528 ; 
   reg __408528_408528;
   reg _408529_408529 ; 
   reg __408529_408529;
   reg _408530_408530 ; 
   reg __408530_408530;
   reg _408531_408531 ; 
   reg __408531_408531;
   reg _408532_408532 ; 
   reg __408532_408532;
   reg _408533_408533 ; 
   reg __408533_408533;
   reg _408534_408534 ; 
   reg __408534_408534;
   reg _408535_408535 ; 
   reg __408535_408535;
   reg _408536_408536 ; 
   reg __408536_408536;
   reg _408537_408537 ; 
   reg __408537_408537;
   reg _408538_408538 ; 
   reg __408538_408538;
   reg _408539_408539 ; 
   reg __408539_408539;
   reg _408540_408540 ; 
   reg __408540_408540;
   reg _408541_408541 ; 
   reg __408541_408541;
   reg _408542_408542 ; 
   reg __408542_408542;
   reg _408543_408543 ; 
   reg __408543_408543;
   reg _408544_408544 ; 
   reg __408544_408544;
   reg _408545_408545 ; 
   reg __408545_408545;
   reg _408546_408546 ; 
   reg __408546_408546;
   reg _408547_408547 ; 
   reg __408547_408547;
   reg _408548_408548 ; 
   reg __408548_408548;
   reg _408549_408549 ; 
   reg __408549_408549;
   reg _408550_408550 ; 
   reg __408550_408550;
   reg _408551_408551 ; 
   reg __408551_408551;
   reg _408552_408552 ; 
   reg __408552_408552;
   reg _408553_408553 ; 
   reg __408553_408553;
   reg _408554_408554 ; 
   reg __408554_408554;
   reg _408555_408555 ; 
   reg __408555_408555;
   reg _408556_408556 ; 
   reg __408556_408556;
   reg _408557_408557 ; 
   reg __408557_408557;
   reg _408558_408558 ; 
   reg __408558_408558;
   reg _408559_408559 ; 
   reg __408559_408559;
   reg _408560_408560 ; 
   reg __408560_408560;
   reg _408561_408561 ; 
   reg __408561_408561;
   reg _408562_408562 ; 
   reg __408562_408562;
   reg _408563_408563 ; 
   reg __408563_408563;
   reg _408564_408564 ; 
   reg __408564_408564;
   reg _408565_408565 ; 
   reg __408565_408565;
   reg _408566_408566 ; 
   reg __408566_408566;
   reg _408567_408567 ; 
   reg __408567_408567;
   reg _408568_408568 ; 
   reg __408568_408568;
   reg _408569_408569 ; 
   reg __408569_408569;
   reg _408570_408570 ; 
   reg __408570_408570;
   reg _408571_408571 ; 
   reg __408571_408571;
   reg _408572_408572 ; 
   reg __408572_408572;
   reg _408573_408573 ; 
   reg __408573_408573;
   reg _408574_408574 ; 
   reg __408574_408574;
   reg _408575_408575 ; 
   reg __408575_408575;
   reg _408576_408576 ; 
   reg __408576_408576;
   reg _408577_408577 ; 
   reg __408577_408577;
   reg _408578_408578 ; 
   reg __408578_408578;
   reg _408579_408579 ; 
   reg __408579_408579;
   reg _408580_408580 ; 
   reg __408580_408580;
   reg _408581_408581 ; 
   reg __408581_408581;
   reg _408582_408582 ; 
   reg __408582_408582;
   reg _408583_408583 ; 
   reg __408583_408583;
   reg _408584_408584 ; 
   reg __408584_408584;
   reg _408585_408585 ; 
   reg __408585_408585;
   reg _408586_408586 ; 
   reg __408586_408586;
   reg _408587_408587 ; 
   reg __408587_408587;
   reg _408588_408588 ; 
   reg __408588_408588;
   reg _408589_408589 ; 
   reg __408589_408589;
   reg _408590_408590 ; 
   reg __408590_408590;
   reg _408591_408591 ; 
   reg __408591_408591;
   reg _408592_408592 ; 
   reg __408592_408592;
   reg _408593_408593 ; 
   reg __408593_408593;
   reg _408594_408594 ; 
   reg __408594_408594;
   reg _408595_408595 ; 
   reg __408595_408595;
   reg _408596_408596 ; 
   reg __408596_408596;
   reg _408597_408597 ; 
   reg __408597_408597;
   reg _408598_408598 ; 
   reg __408598_408598;
   reg _408599_408599 ; 
   reg __408599_408599;
   reg _408600_408600 ; 
   reg __408600_408600;
   reg _408601_408601 ; 
   reg __408601_408601;
   reg _408602_408602 ; 
   reg __408602_408602;
   reg _408603_408603 ; 
   reg __408603_408603;
   reg _408604_408604 ; 
   reg __408604_408604;
   reg _408605_408605 ; 
   reg __408605_408605;
   reg _408606_408606 ; 
   reg __408606_408606;
   reg _408607_408607 ; 
   reg __408607_408607;
   reg _408608_408608 ; 
   reg __408608_408608;
   reg _408609_408609 ; 
   reg __408609_408609;
   reg _408610_408610 ; 
   reg __408610_408610;
   reg _408611_408611 ; 
   reg __408611_408611;
   reg _408612_408612 ; 
   reg __408612_408612;
   reg _408613_408613 ; 
   reg __408613_408613;
   reg _408614_408614 ; 
   reg __408614_408614;
   reg _408615_408615 ; 
   reg __408615_408615;
   reg _408616_408616 ; 
   reg __408616_408616;
   reg _408617_408617 ; 
   reg __408617_408617;
   reg _408618_408618 ; 
   reg __408618_408618;
   reg _408619_408619 ; 
   reg __408619_408619;
   reg _408620_408620 ; 
   reg __408620_408620;
   reg _408621_408621 ; 
   reg __408621_408621;
   reg _408622_408622 ; 
   reg __408622_408622;
   reg _408623_408623 ; 
   reg __408623_408623;
   reg _408624_408624 ; 
   reg __408624_408624;
   reg _408625_408625 ; 
   reg __408625_408625;
   reg _408626_408626 ; 
   reg __408626_408626;
   reg _408627_408627 ; 
   reg __408627_408627;
   reg _408628_408628 ; 
   reg __408628_408628;
   reg _408629_408629 ; 
   reg __408629_408629;
   reg _408630_408630 ; 
   reg __408630_408630;
   reg _408631_408631 ; 
   reg __408631_408631;
   reg _408632_408632 ; 
   reg __408632_408632;
   reg _408633_408633 ; 
   reg __408633_408633;
   reg _408634_408634 ; 
   reg __408634_408634;
   reg _408635_408635 ; 
   reg __408635_408635;
   reg _408636_408636 ; 
   reg __408636_408636;
   reg _408637_408637 ; 
   reg __408637_408637;
   reg _408638_408638 ; 
   reg __408638_408638;
   reg _408639_408639 ; 
   reg __408639_408639;
   reg _408640_408640 ; 
   reg __408640_408640;
   reg _408641_408641 ; 
   reg __408641_408641;
   reg _408642_408642 ; 
   reg __408642_408642;
   reg _408643_408643 ; 
   reg __408643_408643;
   reg _408644_408644 ; 
   reg __408644_408644;
   reg _408645_408645 ; 
   reg __408645_408645;
   reg _408646_408646 ; 
   reg __408646_408646;
   reg _408647_408647 ; 
   reg __408647_408647;
   reg _408648_408648 ; 
   reg __408648_408648;
   reg _408649_408649 ; 
   reg __408649_408649;
   reg _408650_408650 ; 
   reg __408650_408650;
   reg _408651_408651 ; 
   reg __408651_408651;
   reg _408652_408652 ; 
   reg __408652_408652;
   reg _408653_408653 ; 
   reg __408653_408653;
   reg _408654_408654 ; 
   reg __408654_408654;
   reg _408655_408655 ; 
   reg __408655_408655;
   reg _408656_408656 ; 
   reg __408656_408656;
   reg _408657_408657 ; 
   reg __408657_408657;
   reg _408658_408658 ; 
   reg __408658_408658;
   reg _408659_408659 ; 
   reg __408659_408659;
   reg _408660_408660 ; 
   reg __408660_408660;
   reg _408661_408661 ; 
   reg __408661_408661;
   reg _408662_408662 ; 
   reg __408662_408662;
   reg _408663_408663 ; 
   reg __408663_408663;
   reg _408664_408664 ; 
   reg __408664_408664;
   reg _408665_408665 ; 
   reg __408665_408665;
   reg _408666_408666 ; 
   reg __408666_408666;
   reg _408667_408667 ; 
   reg __408667_408667;
   reg _408668_408668 ; 
   reg __408668_408668;
   reg _408669_408669 ; 
   reg __408669_408669;
   reg _408670_408670 ; 
   reg __408670_408670;
   reg _408671_408671 ; 
   reg __408671_408671;
   reg _408672_408672 ; 
   reg __408672_408672;
   reg _408673_408673 ; 
   reg __408673_408673;
   reg _408674_408674 ; 
   reg __408674_408674;
   reg _408675_408675 ; 
   reg __408675_408675;
   reg _408676_408676 ; 
   reg __408676_408676;
   reg _408677_408677 ; 
   reg __408677_408677;
   reg _408678_408678 ; 
   reg __408678_408678;
   reg _408679_408679 ; 
   reg __408679_408679;
   reg _408680_408680 ; 
   reg __408680_408680;
   reg _408681_408681 ; 
   reg __408681_408681;
   reg _408682_408682 ; 
   reg __408682_408682;
   reg _408683_408683 ; 
   reg __408683_408683;
   reg _408684_408684 ; 
   reg __408684_408684;
   reg _408685_408685 ; 
   reg __408685_408685;
   reg _408686_408686 ; 
   reg __408686_408686;
   reg _408687_408687 ; 
   reg __408687_408687;
   reg _408688_408688 ; 
   reg __408688_408688;
   reg _408689_408689 ; 
   reg __408689_408689;
   reg _408690_408690 ; 
   reg __408690_408690;
   reg _408691_408691 ; 
   reg __408691_408691;
   reg _408692_408692 ; 
   reg __408692_408692;
   reg _408693_408693 ; 
   reg __408693_408693;
   reg _408694_408694 ; 
   reg __408694_408694;
   reg _408695_408695 ; 
   reg __408695_408695;
   reg _408696_408696 ; 
   reg __408696_408696;
   reg _408697_408697 ; 
   reg __408697_408697;
   reg _408698_408698 ; 
   reg __408698_408698;
   reg _408699_408699 ; 
   reg __408699_408699;
   reg _408700_408700 ; 
   reg __408700_408700;
   reg _408701_408701 ; 
   reg __408701_408701;
   reg _408702_408702 ; 
   reg __408702_408702;
   reg _408703_408703 ; 
   reg __408703_408703;
   reg _408704_408704 ; 
   reg __408704_408704;
   reg _408705_408705 ; 
   reg __408705_408705;
   reg _408706_408706 ; 
   reg __408706_408706;
   reg _408707_408707 ; 
   reg __408707_408707;
   reg _408708_408708 ; 
   reg __408708_408708;
   reg _408709_408709 ; 
   reg __408709_408709;
   reg _408710_408710 ; 
   reg __408710_408710;
   reg _408711_408711 ; 
   reg __408711_408711;
   reg _408712_408712 ; 
   reg __408712_408712;
   reg _408713_408713 ; 
   reg __408713_408713;
   reg _408714_408714 ; 
   reg __408714_408714;
   reg _408715_408715 ; 
   reg __408715_408715;
   reg _408716_408716 ; 
   reg __408716_408716;
   reg _408717_408717 ; 
   reg __408717_408717;
   reg _408718_408718 ; 
   reg __408718_408718;
   reg _408719_408719 ; 
   reg __408719_408719;
   reg _408720_408720 ; 
   reg __408720_408720;
   reg _408721_408721 ; 
   reg __408721_408721;
   reg _408722_408722 ; 
   reg __408722_408722;
   reg _408723_408723 ; 
   reg __408723_408723;
   reg _408724_408724 ; 
   reg __408724_408724;
   reg _408725_408725 ; 
   reg __408725_408725;
   reg _408726_408726 ; 
   reg __408726_408726;
   reg _408727_408727 ; 
   reg __408727_408727;
   reg _408728_408728 ; 
   reg __408728_408728;
   reg _408729_408729 ; 
   reg __408729_408729;
   reg _408730_408730 ; 
   reg __408730_408730;
   reg _408731_408731 ; 
   reg __408731_408731;
   reg _408732_408732 ; 
   reg __408732_408732;
   reg _408733_408733 ; 
   reg __408733_408733;
   reg _408734_408734 ; 
   reg __408734_408734;
   reg _408735_408735 ; 
   reg __408735_408735;
   reg _408736_408736 ; 
   reg __408736_408736;
   reg _408737_408737 ; 
   reg __408737_408737;
   reg _408738_408738 ; 
   reg __408738_408738;
   reg _408739_408739 ; 
   reg __408739_408739;
   reg _408740_408740 ; 
   reg __408740_408740;
   reg _408741_408741 ; 
   reg __408741_408741;
   reg _408742_408742 ; 
   reg __408742_408742;
   reg _408743_408743 ; 
   reg __408743_408743;
   reg _408744_408744 ; 
   reg __408744_408744;
   reg _408745_408745 ; 
   reg __408745_408745;
   reg _408746_408746 ; 
   reg __408746_408746;
   reg _408747_408747 ; 
   reg __408747_408747;
   reg _408748_408748 ; 
   reg __408748_408748;
   reg _408749_408749 ; 
   reg __408749_408749;
   reg _408750_408750 ; 
   reg __408750_408750;
   reg _408751_408751 ; 
   reg __408751_408751;
   reg _408752_408752 ; 
   reg __408752_408752;
   reg _408753_408753 ; 
   reg __408753_408753;
   reg _408754_408754 ; 
   reg __408754_408754;
   reg _408755_408755 ; 
   reg __408755_408755;
   reg _408756_408756 ; 
   reg __408756_408756;
   reg _408757_408757 ; 
   reg __408757_408757;
   reg _408758_408758 ; 
   reg __408758_408758;
   reg _408759_408759 ; 
   reg __408759_408759;
   reg _408760_408760 ; 
   reg __408760_408760;
   reg _408761_408761 ; 
   reg __408761_408761;
   reg _408762_408762 ; 
   reg __408762_408762;
   reg _408763_408763 ; 
   reg __408763_408763;
   reg _408764_408764 ; 
   reg __408764_408764;
   reg _408765_408765 ; 
   reg __408765_408765;
   reg _408766_408766 ; 
   reg __408766_408766;
   reg _408767_408767 ; 
   reg __408767_408767;
   reg _408768_408768 ; 
   reg __408768_408768;
   reg _408769_408769 ; 
   reg __408769_408769;
   reg _408770_408770 ; 
   reg __408770_408770;
   reg _408771_408771 ; 
   reg __408771_408771;
   reg _408772_408772 ; 
   reg __408772_408772;
   reg _408773_408773 ; 
   reg __408773_408773;
   reg _408774_408774 ; 
   reg __408774_408774;
   reg _408775_408775 ; 
   reg __408775_408775;
   reg _408776_408776 ; 
   reg __408776_408776;
   reg _408777_408777 ; 
   reg __408777_408777;
   reg _408778_408778 ; 
   reg __408778_408778;
   reg _408779_408779 ; 
   reg __408779_408779;
   reg _408780_408780 ; 
   reg __408780_408780;
   reg _408781_408781 ; 
   reg __408781_408781;
   reg _408782_408782 ; 
   reg __408782_408782;
   reg _408783_408783 ; 
   reg __408783_408783;
   reg _408784_408784 ; 
   reg __408784_408784;
   reg _408785_408785 ; 
   reg __408785_408785;
   reg _408786_408786 ; 
   reg __408786_408786;
   reg _408787_408787 ; 
   reg __408787_408787;
   reg _408788_408788 ; 
   reg __408788_408788;
   reg _408789_408789 ; 
   reg __408789_408789;
   reg _408790_408790 ; 
   reg __408790_408790;
   reg _408791_408791 ; 
   reg __408791_408791;
   reg _408792_408792 ; 
   reg __408792_408792;
   reg _408793_408793 ; 
   reg __408793_408793;
   reg _408794_408794 ; 
   reg __408794_408794;
   reg _408795_408795 ; 
   reg __408795_408795;
   reg _408796_408796 ; 
   reg __408796_408796;
   reg _408797_408797 ; 
   reg __408797_408797;
   reg _408798_408798 ; 
   reg __408798_408798;
   reg _408799_408799 ; 
   reg __408799_408799;
   reg _408800_408800 ; 
   reg __408800_408800;
   reg _408801_408801 ; 
   reg __408801_408801;
   reg _408802_408802 ; 
   reg __408802_408802;
   reg _408803_408803 ; 
   reg __408803_408803;
   reg _408804_408804 ; 
   reg __408804_408804;
   reg _408805_408805 ; 
   reg __408805_408805;
   reg _408806_408806 ; 
   reg __408806_408806;
   reg _408807_408807 ; 
   reg __408807_408807;
   reg _408808_408808 ; 
   reg __408808_408808;
   reg _408809_408809 ; 
   reg __408809_408809;
   reg _408810_408810 ; 
   reg __408810_408810;
   reg _408811_408811 ; 
   reg __408811_408811;
   reg _408812_408812 ; 
   reg __408812_408812;
   reg _408813_408813 ; 
   reg __408813_408813;
   reg _408814_408814 ; 
   reg __408814_408814;
   reg _408815_408815 ; 
   reg __408815_408815;
   reg _408816_408816 ; 
   reg __408816_408816;
   reg _408817_408817 ; 
   reg __408817_408817;
   reg _408818_408818 ; 
   reg __408818_408818;
   reg _408819_408819 ; 
   reg __408819_408819;
   reg _408820_408820 ; 
   reg __408820_408820;
   reg _408821_408821 ; 
   reg __408821_408821;
   reg _408822_408822 ; 
   reg __408822_408822;
   reg _408823_408823 ; 
   reg __408823_408823;
   reg _408824_408824 ; 
   reg __408824_408824;
   reg _408825_408825 ; 
   reg __408825_408825;
   reg _408826_408826 ; 
   reg __408826_408826;
   reg _408827_408827 ; 
   reg __408827_408827;
   reg _408828_408828 ; 
   reg __408828_408828;
   reg _408829_408829 ; 
   reg __408829_408829;
   reg _408830_408830 ; 
   reg __408830_408830;
   reg _408831_408831 ; 
   reg __408831_408831;
   reg _408832_408832 ; 
   reg __408832_408832;
   reg _408833_408833 ; 
   reg __408833_408833;
   reg _408834_408834 ; 
   reg __408834_408834;
   reg _408835_408835 ; 
   reg __408835_408835;
   reg _408836_408836 ; 
   reg __408836_408836;
   reg _408837_408837 ; 
   reg __408837_408837;
   reg _408838_408838 ; 
   reg __408838_408838;
   reg _408839_408839 ; 
   reg __408839_408839;
   reg _408840_408840 ; 
   reg __408840_408840;
   reg _408841_408841 ; 
   reg __408841_408841;
   reg _408842_408842 ; 
   reg __408842_408842;
   reg _408843_408843 ; 
   reg __408843_408843;
   reg _408844_408844 ; 
   reg __408844_408844;
   reg _408845_408845 ; 
   reg __408845_408845;
   reg _408846_408846 ; 
   reg __408846_408846;
   reg _408847_408847 ; 
   reg __408847_408847;
   reg _408848_408848 ; 
   reg __408848_408848;
   reg _408849_408849 ; 
   reg __408849_408849;
   reg _408850_408850 ; 
   reg __408850_408850;
   reg _408851_408851 ; 
   reg __408851_408851;
   reg _408852_408852 ; 
   reg __408852_408852;
   reg _408853_408853 ; 
   reg __408853_408853;
   reg _408854_408854 ; 
   reg __408854_408854;
   reg _408855_408855 ; 
   reg __408855_408855;
   reg _408856_408856 ; 
   reg __408856_408856;
   reg _408857_408857 ; 
   reg __408857_408857;
   reg _408858_408858 ; 
   reg __408858_408858;
   reg _408859_408859 ; 
   reg __408859_408859;
   reg _408860_408860 ; 
   reg __408860_408860;
   reg _408861_408861 ; 
   reg __408861_408861;
   reg _408862_408862 ; 
   reg __408862_408862;
   reg _408863_408863 ; 
   reg __408863_408863;
   reg _408864_408864 ; 
   reg __408864_408864;
   reg _408865_408865 ; 
   reg __408865_408865;
   reg _408866_408866 ; 
   reg __408866_408866;
   reg _408867_408867 ; 
   reg __408867_408867;
   reg _408868_408868 ; 
   reg __408868_408868;
   reg _408869_408869 ; 
   reg __408869_408869;
   reg _408870_408870 ; 
   reg __408870_408870;
   reg _408871_408871 ; 
   reg __408871_408871;
   reg _408872_408872 ; 
   reg __408872_408872;
   reg _408873_408873 ; 
   reg __408873_408873;
   reg _408874_408874 ; 
   reg __408874_408874;
   reg _408875_408875 ; 
   reg __408875_408875;
   reg _408876_408876 ; 
   reg __408876_408876;
   reg _408877_408877 ; 
   reg __408877_408877;
   reg _408878_408878 ; 
   reg __408878_408878;
   reg _408879_408879 ; 
   reg __408879_408879;
   reg _408880_408880 ; 
   reg __408880_408880;
   reg _408881_408881 ; 
   reg __408881_408881;
   reg _408882_408882 ; 
   reg __408882_408882;
   reg _408883_408883 ; 
   reg __408883_408883;
   reg _408884_408884 ; 
   reg __408884_408884;
   reg _408885_408885 ; 
   reg __408885_408885;
   reg _408886_408886 ; 
   reg __408886_408886;
   reg _408887_408887 ; 
   reg __408887_408887;
   reg _408888_408888 ; 
   reg __408888_408888;
   reg _408889_408889 ; 
   reg __408889_408889;
   reg _408890_408890 ; 
   reg __408890_408890;
   reg _408891_408891 ; 
   reg __408891_408891;
   reg _408892_408892 ; 
   reg __408892_408892;
   reg _408893_408893 ; 
   reg __408893_408893;
   reg _408894_408894 ; 
   reg __408894_408894;
   reg _408895_408895 ; 
   reg __408895_408895;
   reg _408896_408896 ; 
   reg __408896_408896;
   reg _408897_408897 ; 
   reg __408897_408897;
   reg _408898_408898 ; 
   reg __408898_408898;
   reg _408899_408899 ; 
   reg __408899_408899;
   reg _408900_408900 ; 
   reg __408900_408900;
   reg _408901_408901 ; 
   reg __408901_408901;
   reg _408902_408902 ; 
   reg __408902_408902;
   reg _408903_408903 ; 
   reg __408903_408903;
   reg _408904_408904 ; 
   reg __408904_408904;
   reg _408905_408905 ; 
   reg __408905_408905;
   reg _408906_408906 ; 
   reg __408906_408906;
   reg _408907_408907 ; 
   reg __408907_408907;
   reg _408908_408908 ; 
   reg __408908_408908;
   reg _408909_408909 ; 
   reg __408909_408909;
   reg _408910_408910 ; 
   reg __408910_408910;
   reg _408911_408911 ; 
   reg __408911_408911;
   reg _408912_408912 ; 
   reg __408912_408912;
   reg _408913_408913 ; 
   reg __408913_408913;
   reg _408914_408914 ; 
   reg __408914_408914;
   reg _408915_408915 ; 
   reg __408915_408915;
   reg _408916_408916 ; 
   reg __408916_408916;
   reg _408917_408917 ; 
   reg __408917_408917;
   reg _408918_408918 ; 
   reg __408918_408918;
   reg _408919_408919 ; 
   reg __408919_408919;
   reg _408920_408920 ; 
   reg __408920_408920;
   reg _408921_408921 ; 
   reg __408921_408921;
   reg _408922_408922 ; 
   reg __408922_408922;
   reg _408923_408923 ; 
   reg __408923_408923;
   reg _408924_408924 ; 
   reg __408924_408924;
   reg _408925_408925 ; 
   reg __408925_408925;
   reg _408926_408926 ; 
   reg __408926_408926;
   reg _408927_408927 ; 
   reg __408927_408927;
   reg _408928_408928 ; 
   reg __408928_408928;
   reg _408929_408929 ; 
   reg __408929_408929;
   reg _408930_408930 ; 
   reg __408930_408930;
   reg _408931_408931 ; 
   reg __408931_408931;
   reg _408932_408932 ; 
   reg __408932_408932;
   reg _408933_408933 ; 
   reg __408933_408933;
   reg _408934_408934 ; 
   reg __408934_408934;
   reg _408935_408935 ; 
   reg __408935_408935;
   reg _408936_408936 ; 
   reg __408936_408936;
   reg _408937_408937 ; 
   reg __408937_408937;
   reg _408938_408938 ; 
   reg __408938_408938;
   reg _408939_408939 ; 
   reg __408939_408939;
   reg _408940_408940 ; 
   reg __408940_408940;
   reg _408941_408941 ; 
   reg __408941_408941;
   reg _408942_408942 ; 
   reg __408942_408942;
   reg _408943_408943 ; 
   reg __408943_408943;
   reg _408944_408944 ; 
   reg __408944_408944;
   reg _408945_408945 ; 
   reg __408945_408945;
   reg _408946_408946 ; 
   reg __408946_408946;
   reg _408947_408947 ; 
   reg __408947_408947;
   reg _408948_408948 ; 
   reg __408948_408948;
   reg _408949_408949 ; 
   reg __408949_408949;
   reg _408950_408950 ; 
   reg __408950_408950;
   reg _408951_408951 ; 
   reg __408951_408951;
   reg _408952_408952 ; 
   reg __408952_408952;
   reg _408953_408953 ; 
   reg __408953_408953;
   reg _408954_408954 ; 
   reg __408954_408954;
   reg _408955_408955 ; 
   reg __408955_408955;
   reg _408956_408956 ; 
   reg __408956_408956;
   reg _408957_408957 ; 
   reg __408957_408957;
   reg _408958_408958 ; 
   reg __408958_408958;
   reg _408959_408959 ; 
   reg __408959_408959;
   reg _408960_408960 ; 
   reg __408960_408960;
   reg _408961_408961 ; 
   reg __408961_408961;
   reg _408962_408962 ; 
   reg __408962_408962;
   reg _408963_408963 ; 
   reg __408963_408963;
   reg _408964_408964 ; 
   reg __408964_408964;
   reg _408965_408965 ; 
   reg __408965_408965;
   reg _408966_408966 ; 
   reg __408966_408966;
   reg _408967_408967 ; 
   reg __408967_408967;
   reg _408968_408968 ; 
   reg __408968_408968;
   reg _408969_408969 ; 
   reg __408969_408969;
   reg _408970_408970 ; 
   reg __408970_408970;
   reg _408971_408971 ; 
   reg __408971_408971;
   reg _408972_408972 ; 
   reg __408972_408972;
   reg _408973_408973 ; 
   reg __408973_408973;
   reg _408974_408974 ; 
   reg __408974_408974;
   reg _408975_408975 ; 
   reg __408975_408975;
   reg _408976_408976 ; 
   reg __408976_408976;
   reg _408977_408977 ; 
   reg __408977_408977;
   reg _408978_408978 ; 
   reg __408978_408978;
   reg _408979_408979 ; 
   reg __408979_408979;
   reg _408980_408980 ; 
   reg __408980_408980;
   reg _408981_408981 ; 
   reg __408981_408981;
   reg _408982_408982 ; 
   reg __408982_408982;
   reg _408983_408983 ; 
   reg __408983_408983;
   reg _408984_408984 ; 
   reg __408984_408984;
   reg _408985_408985 ; 
   reg __408985_408985;
   reg _408986_408986 ; 
   reg __408986_408986;
   reg _408987_408987 ; 
   reg __408987_408987;
   reg _408988_408988 ; 
   reg __408988_408988;
   reg _408989_408989 ; 
   reg __408989_408989;
   reg _408990_408990 ; 
   reg __408990_408990;
   reg _408991_408991 ; 
   reg __408991_408991;
   reg _408992_408992 ; 
   reg __408992_408992;
   reg _408993_408993 ; 
   reg __408993_408993;
   reg _408994_408994 ; 
   reg __408994_408994;
   reg _408995_408995 ; 
   reg __408995_408995;
   reg _408996_408996 ; 
   reg __408996_408996;
   reg _408997_408997 ; 
   reg __408997_408997;
   reg _408998_408998 ; 
   reg __408998_408998;
   reg _408999_408999 ; 
   reg __408999_408999;
   reg _409000_409000 ; 
   reg __409000_409000;
   reg _409001_409001 ; 
   reg __409001_409001;
   reg _409002_409002 ; 
   reg __409002_409002;
   reg _409003_409003 ; 
   reg __409003_409003;
   reg _409004_409004 ; 
   reg __409004_409004;
   reg _409005_409005 ; 
   reg __409005_409005;
   reg _409006_409006 ; 
   reg __409006_409006;
   reg _409007_409007 ; 
   reg __409007_409007;
   reg _409008_409008 ; 
   reg __409008_409008;
   reg _409009_409009 ; 
   reg __409009_409009;
   reg _409010_409010 ; 
   reg __409010_409010;
   reg _409011_409011 ; 
   reg __409011_409011;
   reg _409012_409012 ; 
   reg __409012_409012;
   reg _409013_409013 ; 
   reg __409013_409013;
   reg _409014_409014 ; 
   reg __409014_409014;
   reg _409015_409015 ; 
   reg __409015_409015;
   reg _409016_409016 ; 
   reg __409016_409016;
   reg _409017_409017 ; 
   reg __409017_409017;
   reg _409018_409018 ; 
   reg __409018_409018;
   reg _409019_409019 ; 
   reg __409019_409019;
   reg _409020_409020 ; 
   reg __409020_409020;
   reg _409021_409021 ; 
   reg __409021_409021;
   reg _409022_409022 ; 
   reg __409022_409022;
   reg _409023_409023 ; 
   reg __409023_409023;
   reg _409024_409024 ; 
   reg __409024_409024;
   reg _409025_409025 ; 
   reg __409025_409025;
   reg _409026_409026 ; 
   reg __409026_409026;
   reg _409027_409027 ; 
   reg __409027_409027;
   reg _409028_409028 ; 
   reg __409028_409028;
   reg _409029_409029 ; 
   reg __409029_409029;
   reg _409030_409030 ; 
   reg __409030_409030;
   reg _409031_409031 ; 
   reg __409031_409031;
   reg _409032_409032 ; 
   reg __409032_409032;
   reg _409033_409033 ; 
   reg __409033_409033;
   reg _409034_409034 ; 
   reg __409034_409034;
   reg _409035_409035 ; 
   reg __409035_409035;
   reg _409036_409036 ; 
   reg __409036_409036;
   reg _409037_409037 ; 
   reg __409037_409037;
   reg _409038_409038 ; 
   reg __409038_409038;
   reg _409039_409039 ; 
   reg __409039_409039;
   reg _409040_409040 ; 
   reg __409040_409040;
   reg _409041_409041 ; 
   reg __409041_409041;
   reg _409042_409042 ; 
   reg __409042_409042;
   reg _409043_409043 ; 
   reg __409043_409043;
   reg _409044_409044 ; 
   reg __409044_409044;
   reg _409045_409045 ; 
   reg __409045_409045;
   reg _409046_409046 ; 
   reg __409046_409046;
   reg _409047_409047 ; 
   reg __409047_409047;
   reg _409048_409048 ; 
   reg __409048_409048;
   reg _409049_409049 ; 
   reg __409049_409049;
   reg _409050_409050 ; 
   reg __409050_409050;
   reg _409051_409051 ; 
   reg __409051_409051;
   reg _409052_409052 ; 
   reg __409052_409052;
   reg _409053_409053 ; 
   reg __409053_409053;
   reg _409054_409054 ; 
   reg __409054_409054;
   reg _409055_409055 ; 
   reg __409055_409055;
   reg _409056_409056 ; 
   reg __409056_409056;
   reg _409057_409057 ; 
   reg __409057_409057;
   reg _409058_409058 ; 
   reg __409058_409058;
   reg _409059_409059 ; 
   reg __409059_409059;
   reg _409060_409060 ; 
   reg __409060_409060;
   reg _409061_409061 ; 
   reg __409061_409061;
   reg _409062_409062 ; 
   reg __409062_409062;
   reg _409063_409063 ; 
   reg __409063_409063;
   reg _409064_409064 ; 
   reg __409064_409064;
   reg _409065_409065 ; 
   reg __409065_409065;
   reg _409066_409066 ; 
   reg __409066_409066;
   reg _409067_409067 ; 
   reg __409067_409067;
   reg _409068_409068 ; 
   reg __409068_409068;
   reg _409069_409069 ; 
   reg __409069_409069;
   reg _409070_409070 ; 
   reg __409070_409070;
   reg _409071_409071 ; 
   reg __409071_409071;
   reg _409072_409072 ; 
   reg __409072_409072;
   reg _409073_409073 ; 
   reg __409073_409073;
   reg _409074_409074 ; 
   reg __409074_409074;
   reg _409075_409075 ; 
   reg __409075_409075;
   reg _409076_409076 ; 
   reg __409076_409076;
   reg _409077_409077 ; 
   reg __409077_409077;
   reg _409078_409078 ; 
   reg __409078_409078;
   reg _409079_409079 ; 
   reg __409079_409079;
   reg _409080_409080 ; 
   reg __409080_409080;
   reg _409081_409081 ; 
   reg __409081_409081;
   reg _409082_409082 ; 
   reg __409082_409082;
   reg _409083_409083 ; 
   reg __409083_409083;
   reg _409084_409084 ; 
   reg __409084_409084;
   reg _409085_409085 ; 
   reg __409085_409085;
   reg _409086_409086 ; 
   reg __409086_409086;
   reg _409087_409087 ; 
   reg __409087_409087;
   reg _409088_409088 ; 
   reg __409088_409088;
   reg _409089_409089 ; 
   reg __409089_409089;
   reg _409090_409090 ; 
   reg __409090_409090;
   reg _409091_409091 ; 
   reg __409091_409091;
   reg _409092_409092 ; 
   reg __409092_409092;
   reg _409093_409093 ; 
   reg __409093_409093;
   reg _409094_409094 ; 
   reg __409094_409094;
   reg _409095_409095 ; 
   reg __409095_409095;
   reg _409096_409096 ; 
   reg __409096_409096;
   reg _409097_409097 ; 
   reg __409097_409097;
   reg _409098_409098 ; 
   reg __409098_409098;
   reg _409099_409099 ; 
   reg __409099_409099;
   reg _409100_409100 ; 
   reg __409100_409100;
   reg _409101_409101 ; 
   reg __409101_409101;
   reg _409102_409102 ; 
   reg __409102_409102;
   reg _409103_409103 ; 
   reg __409103_409103;
   reg _409104_409104 ; 
   reg __409104_409104;
   reg _409105_409105 ; 
   reg __409105_409105;
   reg _409106_409106 ; 
   reg __409106_409106;
   reg _409107_409107 ; 
   reg __409107_409107;
   reg _409108_409108 ; 
   reg __409108_409108;
   reg _409109_409109 ; 
   reg __409109_409109;
   reg _409110_409110 ; 
   reg __409110_409110;
   reg _409111_409111 ; 
   reg __409111_409111;
   reg _409112_409112 ; 
   reg __409112_409112;
   reg _409113_409113 ; 
   reg __409113_409113;
   reg _409114_409114 ; 
   reg __409114_409114;
   reg _409115_409115 ; 
   reg __409115_409115;
   reg _409116_409116 ; 
   reg __409116_409116;
   reg _409117_409117 ; 
   reg __409117_409117;
   reg _409118_409118 ; 
   reg __409118_409118;
   reg _409119_409119 ; 
   reg __409119_409119;
   reg _409120_409120 ; 
   reg __409120_409120;
   reg _409121_409121 ; 
   reg __409121_409121;
   reg _409122_409122 ; 
   reg __409122_409122;
   reg _409123_409123 ; 
   reg __409123_409123;
   reg _409124_409124 ; 
   reg __409124_409124;
   reg _409125_409125 ; 
   reg __409125_409125;
   reg _409126_409126 ; 
   reg __409126_409126;
   reg _409127_409127 ; 
   reg __409127_409127;
   reg _409128_409128 ; 
   reg __409128_409128;
   reg _409129_409129 ; 
   reg __409129_409129;
   reg _409130_409130 ; 
   reg __409130_409130;
   reg _409131_409131 ; 
   reg __409131_409131;
   reg _409132_409132 ; 
   reg __409132_409132;
   reg _409133_409133 ; 
   reg __409133_409133;
   reg _409134_409134 ; 
   reg __409134_409134;
   reg _409135_409135 ; 
   reg __409135_409135;
   reg _409136_409136 ; 
   reg __409136_409136;
   reg _409137_409137 ; 
   reg __409137_409137;
   reg _409138_409138 ; 
   reg __409138_409138;
   reg _409139_409139 ; 
   reg __409139_409139;
   reg _409140_409140 ; 
   reg __409140_409140;
   reg _409141_409141 ; 
   reg __409141_409141;
   reg _409142_409142 ; 
   reg __409142_409142;
   reg _409143_409143 ; 
   reg __409143_409143;
   reg _409144_409144 ; 
   reg __409144_409144;
   reg _409145_409145 ; 
   reg __409145_409145;
   reg _409146_409146 ; 
   reg __409146_409146;
   reg _409147_409147 ; 
   reg __409147_409147;
   reg _409148_409148 ; 
   reg __409148_409148;
   reg _409149_409149 ; 
   reg __409149_409149;
   reg _409150_409150 ; 
   reg __409150_409150;
   reg _409151_409151 ; 
   reg __409151_409151;
   reg _409152_409152 ; 
   reg __409152_409152;
   reg _409153_409153 ; 
   reg __409153_409153;
   reg _409154_409154 ; 
   reg __409154_409154;
   reg _409155_409155 ; 
   reg __409155_409155;
   reg _409156_409156 ; 
   reg __409156_409156;
   reg _409157_409157 ; 
   reg __409157_409157;
   reg _409158_409158 ; 
   reg __409158_409158;
   reg _409159_409159 ; 
   reg __409159_409159;
   reg _409160_409160 ; 
   reg __409160_409160;
   reg _409161_409161 ; 
   reg __409161_409161;
   reg _409162_409162 ; 
   reg __409162_409162;
   reg _409163_409163 ; 
   reg __409163_409163;
   reg _409164_409164 ; 
   reg __409164_409164;
   reg _409165_409165 ; 
   reg __409165_409165;
   reg _409166_409166 ; 
   reg __409166_409166;
   reg _409167_409167 ; 
   reg __409167_409167;
   reg _409168_409168 ; 
   reg __409168_409168;
   reg _409169_409169 ; 
   reg __409169_409169;
   reg _409170_409170 ; 
   reg __409170_409170;
   reg _409171_409171 ; 
   reg __409171_409171;
   reg _409172_409172 ; 
   reg __409172_409172;
   reg _409173_409173 ; 
   reg __409173_409173;
   reg _409174_409174 ; 
   reg __409174_409174;
   reg _409175_409175 ; 
   reg __409175_409175;
   reg _409176_409176 ; 
   reg __409176_409176;
   reg _409177_409177 ; 
   reg __409177_409177;
   reg _409178_409178 ; 
   reg __409178_409178;
   reg _409179_409179 ; 
   reg __409179_409179;
   reg _409180_409180 ; 
   reg __409180_409180;
   reg _409181_409181 ; 
   reg __409181_409181;
   reg _409182_409182 ; 
   reg __409182_409182;
   reg _409183_409183 ; 
   reg __409183_409183;
   reg _409184_409184 ; 
   reg __409184_409184;
   reg _409185_409185 ; 
   reg __409185_409185;
   reg _409186_409186 ; 
   reg __409186_409186;
   reg _409187_409187 ; 
   reg __409187_409187;
   reg _409188_409188 ; 
   reg __409188_409188;
   reg _409189_409189 ; 
   reg __409189_409189;
   reg _409190_409190 ; 
   reg __409190_409190;
   reg _409191_409191 ; 
   reg __409191_409191;
   reg _409192_409192 ; 
   reg __409192_409192;
   reg _409193_409193 ; 
   reg __409193_409193;
   reg _409194_409194 ; 
   reg __409194_409194;
   reg _409195_409195 ; 
   reg __409195_409195;
   reg _409196_409196 ; 
   reg __409196_409196;
   reg _409197_409197 ; 
   reg __409197_409197;
   reg _409198_409198 ; 
   reg __409198_409198;
   reg _409199_409199 ; 
   reg __409199_409199;
   reg _409200_409200 ; 
   reg __409200_409200;
   reg _409201_409201 ; 
   reg __409201_409201;
   reg _409202_409202 ; 
   reg __409202_409202;
   reg _409203_409203 ; 
   reg __409203_409203;
   reg _409204_409204 ; 
   reg __409204_409204;
   reg _409205_409205 ; 
   reg __409205_409205;
   reg _409206_409206 ; 
   reg __409206_409206;
   reg _409207_409207 ; 
   reg __409207_409207;
   reg _409208_409208 ; 
   reg __409208_409208;
   reg _409209_409209 ; 
   reg __409209_409209;
   reg _409210_409210 ; 
   reg __409210_409210;
   reg _409211_409211 ; 
   reg __409211_409211;
   reg _409212_409212 ; 
   reg __409212_409212;
   reg _409213_409213 ; 
   reg __409213_409213;
   reg _409214_409214 ; 
   reg __409214_409214;
   reg _409215_409215 ; 
   reg __409215_409215;
   reg _409216_409216 ; 
   reg __409216_409216;
   reg _409217_409217 ; 
   reg __409217_409217;
   reg _409218_409218 ; 
   reg __409218_409218;
   reg _409219_409219 ; 
   reg __409219_409219;
   reg _409220_409220 ; 
   reg __409220_409220;
   reg _409221_409221 ; 
   reg __409221_409221;
   reg _409222_409222 ; 
   reg __409222_409222;
   reg _409223_409223 ; 
   reg __409223_409223;
   reg _409224_409224 ; 
   reg __409224_409224;
   reg _409225_409225 ; 
   reg __409225_409225;
   reg _409226_409226 ; 
   reg __409226_409226;
   reg _409227_409227 ; 
   reg __409227_409227;
   reg _409228_409228 ; 
   reg __409228_409228;
   reg _409229_409229 ; 
   reg __409229_409229;
   reg _409230_409230 ; 
   reg __409230_409230;
   reg _409231_409231 ; 
   reg __409231_409231;
   reg _409232_409232 ; 
   reg __409232_409232;
   reg _409233_409233 ; 
   reg __409233_409233;
   reg _409234_409234 ; 
   reg __409234_409234;
   reg _409235_409235 ; 
   reg __409235_409235;
   reg _409236_409236 ; 
   reg __409236_409236;
   reg _409237_409237 ; 
   reg __409237_409237;
   reg _409238_409238 ; 
   reg __409238_409238;
   reg _409239_409239 ; 
   reg __409239_409239;
   reg _409240_409240 ; 
   reg __409240_409240;
   reg _409241_409241 ; 
   reg __409241_409241;
   reg _409242_409242 ; 
   reg __409242_409242;
   reg _409243_409243 ; 
   reg __409243_409243;
   reg _409244_409244 ; 
   reg __409244_409244;
   reg _409245_409245 ; 
   reg __409245_409245;
   reg _409246_409246 ; 
   reg __409246_409246;
   reg _409247_409247 ; 
   reg __409247_409247;
   reg _409248_409248 ; 
   reg __409248_409248;
   reg _409249_409249 ; 
   reg __409249_409249;
   reg _409250_409250 ; 
   reg __409250_409250;
   reg _409251_409251 ; 
   reg __409251_409251;
   reg _409252_409252 ; 
   reg __409252_409252;
   reg _409253_409253 ; 
   reg __409253_409253;
   reg _409254_409254 ; 
   reg __409254_409254;
   reg _409255_409255 ; 
   reg __409255_409255;
   reg _409256_409256 ; 
   reg __409256_409256;
   reg _409257_409257 ; 
   reg __409257_409257;
   reg _409258_409258 ; 
   reg __409258_409258;
   reg _409259_409259 ; 
   reg __409259_409259;
   reg _409260_409260 ; 
   reg __409260_409260;
   reg _409261_409261 ; 
   reg __409261_409261;
   reg _409262_409262 ; 
   reg __409262_409262;
   reg _409263_409263 ; 
   reg __409263_409263;
   reg _409264_409264 ; 
   reg __409264_409264;
   reg _409265_409265 ; 
   reg __409265_409265;
   reg _409266_409266 ; 
   reg __409266_409266;
   reg _409267_409267 ; 
   reg __409267_409267;
   reg _409268_409268 ; 
   reg __409268_409268;
   reg _409269_409269 ; 
   reg __409269_409269;
   reg _409270_409270 ; 
   reg __409270_409270;
   reg _409271_409271 ; 
   reg __409271_409271;
   reg _409272_409272 ; 
   reg __409272_409272;
   reg _409273_409273 ; 
   reg __409273_409273;
   reg _409274_409274 ; 
   reg __409274_409274;
   reg _409275_409275 ; 
   reg __409275_409275;
   reg _409276_409276 ; 
   reg __409276_409276;
   reg _409277_409277 ; 
   reg __409277_409277;
   reg _409278_409278 ; 
   reg __409278_409278;
   reg _409279_409279 ; 
   reg __409279_409279;
   reg _409280_409280 ; 
   reg __409280_409280;
   reg _409281_409281 ; 
   reg __409281_409281;
   reg _409282_409282 ; 
   reg __409282_409282;
   reg _409283_409283 ; 
   reg __409283_409283;
   reg _409284_409284 ; 
   reg __409284_409284;
   reg _409285_409285 ; 
   reg __409285_409285;
   reg _409286_409286 ; 
   reg __409286_409286;
   reg _409287_409287 ; 
   reg __409287_409287;
   reg _409288_409288 ; 
   reg __409288_409288;
   reg _409289_409289 ; 
   reg __409289_409289;
   reg _409290_409290 ; 
   reg __409290_409290;
   reg _409291_409291 ; 
   reg __409291_409291;
   reg _409292_409292 ; 
   reg __409292_409292;
   reg _409293_409293 ; 
   reg __409293_409293;
   reg _409294_409294 ; 
   reg __409294_409294;
   reg _409295_409295 ; 
   reg __409295_409295;
   reg _409296_409296 ; 
   reg __409296_409296;
   reg _409297_409297 ; 
   reg __409297_409297;
   reg _409298_409298 ; 
   reg __409298_409298;
   reg _409299_409299 ; 
   reg __409299_409299;
   reg _409300_409300 ; 
   reg __409300_409300;
   reg _409301_409301 ; 
   reg __409301_409301;
   reg _409302_409302 ; 
   reg __409302_409302;
   reg _409303_409303 ; 
   reg __409303_409303;
   reg _409304_409304 ; 
   reg __409304_409304;
   reg _409305_409305 ; 
   reg __409305_409305;
   reg _409306_409306 ; 
   reg __409306_409306;
   reg _409307_409307 ; 
   reg __409307_409307;
   reg _409308_409308 ; 
   reg __409308_409308;
   reg _409309_409309 ; 
   reg __409309_409309;
   reg _409310_409310 ; 
   reg __409310_409310;
   reg _409311_409311 ; 
   reg __409311_409311;
   reg _409312_409312 ; 
   reg __409312_409312;
   reg _409313_409313 ; 
   reg __409313_409313;
   reg _409314_409314 ; 
   reg __409314_409314;
   reg _409315_409315 ; 
   reg __409315_409315;
   reg _409316_409316 ; 
   reg __409316_409316;
   reg _409317_409317 ; 
   reg __409317_409317;
   reg _409318_409318 ; 
   reg __409318_409318;
   reg _409319_409319 ; 
   reg __409319_409319;
   reg _409320_409320 ; 
   reg __409320_409320;
   reg _409321_409321 ; 
   reg __409321_409321;
   reg _409322_409322 ; 
   reg __409322_409322;
   reg _409323_409323 ; 
   reg __409323_409323;
   reg _409324_409324 ; 
   reg __409324_409324;
   reg _409325_409325 ; 
   reg __409325_409325;
   reg _409326_409326 ; 
   reg __409326_409326;
   reg _409327_409327 ; 
   reg __409327_409327;
   reg _409328_409328 ; 
   reg __409328_409328;
   reg _409329_409329 ; 
   reg __409329_409329;
   reg _409330_409330 ; 
   reg __409330_409330;
   reg _409331_409331 ; 
   reg __409331_409331;
   reg _409332_409332 ; 
   reg __409332_409332;
   reg _409333_409333 ; 
   reg __409333_409333;
   reg _409334_409334 ; 
   reg __409334_409334;
   reg _409335_409335 ; 
   reg __409335_409335;
   reg _409336_409336 ; 
   reg __409336_409336;
   reg _409337_409337 ; 
   reg __409337_409337;
   reg _409338_409338 ; 
   reg __409338_409338;
   reg _409339_409339 ; 
   reg __409339_409339;
   reg _409340_409340 ; 
   reg __409340_409340;
   reg _409341_409341 ; 
   reg __409341_409341;
   reg _409342_409342 ; 
   reg __409342_409342;
   reg _409343_409343 ; 
   reg __409343_409343;
   reg _409344_409344 ; 
   reg __409344_409344;
   reg _409345_409345 ; 
   reg __409345_409345;
   reg _409346_409346 ; 
   reg __409346_409346;
   reg _409347_409347 ; 
   reg __409347_409347;
   reg _409348_409348 ; 
   reg __409348_409348;
   reg _409349_409349 ; 
   reg __409349_409349;
   reg _409350_409350 ; 
   reg __409350_409350;
   reg _409351_409351 ; 
   reg __409351_409351;
   reg _409352_409352 ; 
   reg __409352_409352;
   reg _409353_409353 ; 
   reg __409353_409353;
   reg _409354_409354 ; 
   reg __409354_409354;
   reg _409355_409355 ; 
   reg __409355_409355;
   reg _409356_409356 ; 
   reg __409356_409356;
   reg _409357_409357 ; 
   reg __409357_409357;
   reg _409358_409358 ; 
   reg __409358_409358;
   reg _409359_409359 ; 
   reg __409359_409359;
   reg _409360_409360 ; 
   reg __409360_409360;
   reg _409361_409361 ; 
   reg __409361_409361;
   reg _409362_409362 ; 
   reg __409362_409362;
   reg _409363_409363 ; 
   reg __409363_409363;
   reg _409364_409364 ; 
   reg __409364_409364;
   reg _409365_409365 ; 
   reg __409365_409365;
   reg _409366_409366 ; 
   reg __409366_409366;
   reg _409367_409367 ; 
   reg __409367_409367;
   reg _409368_409368 ; 
   reg __409368_409368;
   reg _409369_409369 ; 
   reg __409369_409369;
   reg _409370_409370 ; 
   reg __409370_409370;
   reg _409371_409371 ; 
   reg __409371_409371;
   reg _409372_409372 ; 
   reg __409372_409372;
   reg _409373_409373 ; 
   reg __409373_409373;
   reg _409374_409374 ; 
   reg __409374_409374;
   reg _409375_409375 ; 
   reg __409375_409375;
   reg _409376_409376 ; 
   reg __409376_409376;
   reg _409377_409377 ; 
   reg __409377_409377;
   reg _409378_409378 ; 
   reg __409378_409378;
   reg _409379_409379 ; 
   reg __409379_409379;
   reg _409380_409380 ; 
   reg __409380_409380;
   reg _409381_409381 ; 
   reg __409381_409381;
   reg _409382_409382 ; 
   reg __409382_409382;
   reg _409383_409383 ; 
   reg __409383_409383;
   reg _409384_409384 ; 
   reg __409384_409384;
   reg _409385_409385 ; 
   reg __409385_409385;
   reg _409386_409386 ; 
   reg __409386_409386;
   reg _409387_409387 ; 
   reg __409387_409387;
   reg _409388_409388 ; 
   reg __409388_409388;
   reg _409389_409389 ; 
   reg __409389_409389;
   reg _409390_409390 ; 
   reg __409390_409390;
   reg _409391_409391 ; 
   reg __409391_409391;
   reg _409392_409392 ; 
   reg __409392_409392;
   reg _409393_409393 ; 
   reg __409393_409393;
   reg _409394_409394 ; 
   reg __409394_409394;
   reg _409395_409395 ; 
   reg __409395_409395;
   reg _409396_409396 ; 
   reg __409396_409396;
   reg _409397_409397 ; 
   reg __409397_409397;
   reg _409398_409398 ; 
   reg __409398_409398;
   reg _409399_409399 ; 
   reg __409399_409399;
   reg _409400_409400 ; 
   reg __409400_409400;
   reg _409401_409401 ; 
   reg __409401_409401;
   reg _409402_409402 ; 
   reg __409402_409402;
   reg _409403_409403 ; 
   reg __409403_409403;
   reg _409404_409404 ; 
   reg __409404_409404;
   reg _409405_409405 ; 
   reg __409405_409405;
   reg _409406_409406 ; 
   reg __409406_409406;
   reg _409407_409407 ; 
   reg __409407_409407;
   reg _409408_409408 ; 
   reg __409408_409408;
   reg _409409_409409 ; 
   reg __409409_409409;
   reg _409410_409410 ; 
   reg __409410_409410;
   reg _409411_409411 ; 
   reg __409411_409411;
   reg _409412_409412 ; 
   reg __409412_409412;
   reg _409413_409413 ; 
   reg __409413_409413;
   reg _409414_409414 ; 
   reg __409414_409414;
   reg _409415_409415 ; 
   reg __409415_409415;
   reg _409416_409416 ; 
   reg __409416_409416;
   reg _409417_409417 ; 
   reg __409417_409417;
   reg _409418_409418 ; 
   reg __409418_409418;
   reg _409419_409419 ; 
   reg __409419_409419;
   reg _409420_409420 ; 
   reg __409420_409420;
   reg _409421_409421 ; 
   reg __409421_409421;
   reg _409422_409422 ; 
   reg __409422_409422;
   reg _409423_409423 ; 
   reg __409423_409423;
   reg _409424_409424 ; 
   reg __409424_409424;
   reg _409425_409425 ; 
   reg __409425_409425;
   reg _409426_409426 ; 
   reg __409426_409426;
   reg _409427_409427 ; 
   reg __409427_409427;
   reg _409428_409428 ; 
   reg __409428_409428;
   reg _409429_409429 ; 
   reg __409429_409429;
   reg _409430_409430 ; 
   reg __409430_409430;
   reg _409431_409431 ; 
   reg __409431_409431;
   reg _409432_409432 ; 
   reg __409432_409432;
   reg _409433_409433 ; 
   reg __409433_409433;
   reg _409434_409434 ; 
   reg __409434_409434;
   reg _409435_409435 ; 
   reg __409435_409435;
   reg _409436_409436 ; 
   reg __409436_409436;
   reg _409437_409437 ; 
   reg __409437_409437;
   reg _409438_409438 ; 
   reg __409438_409438;
   reg _409439_409439 ; 
   reg __409439_409439;
   reg _409440_409440 ; 
   reg __409440_409440;
   reg _409441_409441 ; 
   reg __409441_409441;
   reg _409442_409442 ; 
   reg __409442_409442;
   reg _409443_409443 ; 
   reg __409443_409443;
   reg _409444_409444 ; 
   reg __409444_409444;
   reg _409445_409445 ; 
   reg __409445_409445;
   reg _409446_409446 ; 
   reg __409446_409446;
   reg _409447_409447 ; 
   reg __409447_409447;
   reg _409448_409448 ; 
   reg __409448_409448;
   reg _409449_409449 ; 
   reg __409449_409449;
   reg _409450_409450 ; 
   reg __409450_409450;
   reg _409451_409451 ; 
   reg __409451_409451;
   reg _409452_409452 ; 
   reg __409452_409452;
   reg _409453_409453 ; 
   reg __409453_409453;
   reg _409454_409454 ; 
   reg __409454_409454;
   reg _409455_409455 ; 
   reg __409455_409455;
   reg _409456_409456 ; 
   reg __409456_409456;
   reg _409457_409457 ; 
   reg __409457_409457;
   reg _409458_409458 ; 
   reg __409458_409458;
   reg _409459_409459 ; 
   reg __409459_409459;
   reg _409460_409460 ; 
   reg __409460_409460;
   reg _409461_409461 ; 
   reg __409461_409461;
   reg _409462_409462 ; 
   reg __409462_409462;
   reg _409463_409463 ; 
   reg __409463_409463;
   reg _409464_409464 ; 
   reg __409464_409464;
   reg _409465_409465 ; 
   reg __409465_409465;
   reg _409466_409466 ; 
   reg __409466_409466;
   reg _409467_409467 ; 
   reg __409467_409467;
   reg _409468_409468 ; 
   reg __409468_409468;
   reg _409469_409469 ; 
   reg __409469_409469;
   reg _409470_409470 ; 
   reg __409470_409470;
   reg _409471_409471 ; 
   reg __409471_409471;
   reg _409472_409472 ; 
   reg __409472_409472;
   reg _409473_409473 ; 
   reg __409473_409473;
   reg _409474_409474 ; 
   reg __409474_409474;
   reg _409475_409475 ; 
   reg __409475_409475;
   reg _409476_409476 ; 
   reg __409476_409476;
   reg _409477_409477 ; 
   reg __409477_409477;
   reg _409478_409478 ; 
   reg __409478_409478;
   reg _409479_409479 ; 
   reg __409479_409479;
   reg _409480_409480 ; 
   reg __409480_409480;
   reg _409481_409481 ; 
   reg __409481_409481;
   reg _409482_409482 ; 
   reg __409482_409482;
   reg _409483_409483 ; 
   reg __409483_409483;
   reg _409484_409484 ; 
   reg __409484_409484;
   reg _409485_409485 ; 
   reg __409485_409485;
   reg _409486_409486 ; 
   reg __409486_409486;
   reg _409487_409487 ; 
   reg __409487_409487;
   reg _409488_409488 ; 
   reg __409488_409488;
   reg _409489_409489 ; 
   reg __409489_409489;
   reg _409490_409490 ; 
   reg __409490_409490;
   reg _409491_409491 ; 
   reg __409491_409491;
   reg _409492_409492 ; 
   reg __409492_409492;
   reg _409493_409493 ; 
   reg __409493_409493;
   reg _409494_409494 ; 
   reg __409494_409494;
   reg _409495_409495 ; 
   reg __409495_409495;
   reg _409496_409496 ; 
   reg __409496_409496;
   reg _409497_409497 ; 
   reg __409497_409497;
   reg _409498_409498 ; 
   reg __409498_409498;
   reg _409499_409499 ; 
   reg __409499_409499;
   reg _409500_409500 ; 
   reg __409500_409500;
   reg _409501_409501 ; 
   reg __409501_409501;
   reg _409502_409502 ; 
   reg __409502_409502;
   reg _409503_409503 ; 
   reg __409503_409503;
   reg _409504_409504 ; 
   reg __409504_409504;
   reg _409505_409505 ; 
   reg __409505_409505;
   reg _409506_409506 ; 
   reg __409506_409506;
   reg _409507_409507 ; 
   reg __409507_409507;
   reg _409508_409508 ; 
   reg __409508_409508;
   reg _409509_409509 ; 
   reg __409509_409509;
   reg _409510_409510 ; 
   reg __409510_409510;
   reg _409511_409511 ; 
   reg __409511_409511;
   reg _409512_409512 ; 
   reg __409512_409512;
   reg _409513_409513 ; 
   reg __409513_409513;
   reg _409514_409514 ; 
   reg __409514_409514;
   reg _409515_409515 ; 
   reg __409515_409515;
   reg _409516_409516 ; 
   reg __409516_409516;
   reg _409517_409517 ; 
   reg __409517_409517;
   reg _409518_409518 ; 
   reg __409518_409518;
   reg _409519_409519 ; 
   reg __409519_409519;
   reg _409520_409520 ; 
   reg __409520_409520;
   reg _409521_409521 ; 
   reg __409521_409521;
   reg _409522_409522 ; 
   reg __409522_409522;
   reg _409523_409523 ; 
   reg __409523_409523;
   reg _409524_409524 ; 
   reg __409524_409524;
   reg _409525_409525 ; 
   reg __409525_409525;
   reg _409526_409526 ; 
   reg __409526_409526;
   reg _409527_409527 ; 
   reg __409527_409527;
   reg _409528_409528 ; 
   reg __409528_409528;
   reg _409529_409529 ; 
   reg __409529_409529;
   reg _409530_409530 ; 
   reg __409530_409530;
   reg _409531_409531 ; 
   reg __409531_409531;
   reg _409532_409532 ; 
   reg __409532_409532;
   reg _409533_409533 ; 
   reg __409533_409533;
   reg _409534_409534 ; 
   reg __409534_409534;
   reg _409535_409535 ; 
   reg __409535_409535;
   reg _409536_409536 ; 
   reg __409536_409536;
   reg _409537_409537 ; 
   reg __409537_409537;
   reg _409538_409538 ; 
   reg __409538_409538;
   reg _409539_409539 ; 
   reg __409539_409539;
   reg _409540_409540 ; 
   reg __409540_409540;
   reg _409541_409541 ; 
   reg __409541_409541;
   reg _409542_409542 ; 
   reg __409542_409542;
   reg _409543_409543 ; 
   reg __409543_409543;
   reg _409544_409544 ; 
   reg __409544_409544;
   reg _409545_409545 ; 
   reg __409545_409545;
   reg _409546_409546 ; 
   reg __409546_409546;
   reg _409547_409547 ; 
   reg __409547_409547;
   reg _409548_409548 ; 
   reg __409548_409548;
   reg _409549_409549 ; 
   reg __409549_409549;
   reg _409550_409550 ; 
   reg __409550_409550;
   reg _409551_409551 ; 
   reg __409551_409551;
   reg _409552_409552 ; 
   reg __409552_409552;
   reg _409553_409553 ; 
   reg __409553_409553;
   reg _409554_409554 ; 
   reg __409554_409554;
   reg _409555_409555 ; 
   reg __409555_409555;
   reg _409556_409556 ; 
   reg __409556_409556;
   reg _409557_409557 ; 
   reg __409557_409557;
   reg _409558_409558 ; 
   reg __409558_409558;
   reg _409559_409559 ; 
   reg __409559_409559;
   reg _409560_409560 ; 
   reg __409560_409560;
   reg _409561_409561 ; 
   reg __409561_409561;
   reg _409562_409562 ; 
   reg __409562_409562;
   reg _409563_409563 ; 
   reg __409563_409563;
   reg _409564_409564 ; 
   reg __409564_409564;
   reg _409565_409565 ; 
   reg __409565_409565;
   reg _409566_409566 ; 
   reg __409566_409566;
   reg _409567_409567 ; 
   reg __409567_409567;
   reg _409568_409568 ; 
   reg __409568_409568;
   reg _409569_409569 ; 
   reg __409569_409569;
   reg _409570_409570 ; 
   reg __409570_409570;
   reg _409571_409571 ; 
   reg __409571_409571;
   reg _409572_409572 ; 
   reg __409572_409572;
   reg _409573_409573 ; 
   reg __409573_409573;
   reg _409574_409574 ; 
   reg __409574_409574;
   reg _409575_409575 ; 
   reg __409575_409575;
   reg _409576_409576 ; 
   reg __409576_409576;
   reg _409577_409577 ; 
   reg __409577_409577;
   reg _409578_409578 ; 
   reg __409578_409578;
   reg _409579_409579 ; 
   reg __409579_409579;
   reg _409580_409580 ; 
   reg __409580_409580;
   reg _409581_409581 ; 
   reg __409581_409581;
   reg _409582_409582 ; 
   reg __409582_409582;
   reg _409583_409583 ; 
   reg __409583_409583;
   reg _409584_409584 ; 
   reg __409584_409584;
   reg _409585_409585 ; 
   reg __409585_409585;
   reg _409586_409586 ; 
   reg __409586_409586;
   reg _409587_409587 ; 
   reg __409587_409587;
   reg _409588_409588 ; 
   reg __409588_409588;
   reg _409589_409589 ; 
   reg __409589_409589;
   reg _409590_409590 ; 
   reg __409590_409590;
   reg _409591_409591 ; 
   reg __409591_409591;
   reg _409592_409592 ; 
   reg __409592_409592;
   reg _409593_409593 ; 
   reg __409593_409593;
   reg _409594_409594 ; 
   reg __409594_409594;
   reg _409595_409595 ; 
   reg __409595_409595;
   reg _409596_409596 ; 
   reg __409596_409596;
   reg _409597_409597 ; 
   reg __409597_409597;
   reg _409598_409598 ; 
   reg __409598_409598;
   reg _409599_409599 ; 
   reg __409599_409599;
   reg _409600_409600 ; 
   reg __409600_409600;
   reg _409601_409601 ; 
   reg __409601_409601;
   reg _409602_409602 ; 
   reg __409602_409602;
   reg _409603_409603 ; 
   reg __409603_409603;
   reg _409604_409604 ; 
   reg __409604_409604;
   reg _409605_409605 ; 
   reg __409605_409605;
   reg _409606_409606 ; 
   reg __409606_409606;
   reg _409607_409607 ; 
   reg __409607_409607;
   reg _409608_409608 ; 
   reg __409608_409608;
   reg _409609_409609 ; 
   reg __409609_409609;
   reg _409610_409610 ; 
   reg __409610_409610;
   reg _409611_409611 ; 
   reg __409611_409611;
   reg _409612_409612 ; 
   reg __409612_409612;
   reg _409613_409613 ; 
   reg __409613_409613;
   reg _409614_409614 ; 
   reg __409614_409614;
   reg _409615_409615 ; 
   reg __409615_409615;
   reg _409616_409616 ; 
   reg __409616_409616;
   reg _409617_409617 ; 
   reg __409617_409617;
   reg _409618_409618 ; 
   reg __409618_409618;
   reg _409619_409619 ; 
   reg __409619_409619;
   reg _409620_409620 ; 
   reg __409620_409620;
   reg _409621_409621 ; 
   reg __409621_409621;
   reg _409622_409622 ; 
   reg __409622_409622;
   reg _409623_409623 ; 
   reg __409623_409623;
   reg _409624_409624 ; 
   reg __409624_409624;
   reg _409625_409625 ; 
   reg __409625_409625;
   reg _409626_409626 ; 
   reg __409626_409626;
   reg _409627_409627 ; 
   reg __409627_409627;
   reg _409628_409628 ; 
   reg __409628_409628;
   reg _409629_409629 ; 
   reg __409629_409629;
   reg _409630_409630 ; 
   reg __409630_409630;
   reg _409631_409631 ; 
   reg __409631_409631;
   reg _409632_409632 ; 
   reg __409632_409632;
   reg _409633_409633 ; 
   reg __409633_409633;
   reg _409634_409634 ; 
   reg __409634_409634;
   reg _409635_409635 ; 
   reg __409635_409635;
   reg _409636_409636 ; 
   reg __409636_409636;
   reg _409637_409637 ; 
   reg __409637_409637;
   reg _409638_409638 ; 
   reg __409638_409638;
   reg _409639_409639 ; 
   reg __409639_409639;
   reg _409640_409640 ; 
   reg __409640_409640;
   reg _409641_409641 ; 
   reg __409641_409641;
   reg _409642_409642 ; 
   reg __409642_409642;
   reg _409643_409643 ; 
   reg __409643_409643;
   reg _409644_409644 ; 
   reg __409644_409644;
   reg _409645_409645 ; 
   reg __409645_409645;
   reg _409646_409646 ; 
   reg __409646_409646;
   reg _409647_409647 ; 
   reg __409647_409647;
   reg _409648_409648 ; 
   reg __409648_409648;
   reg _409649_409649 ; 
   reg __409649_409649;
   reg _409650_409650 ; 
   reg __409650_409650;
   reg _409651_409651 ; 
   reg __409651_409651;
   reg _409652_409652 ; 
   reg __409652_409652;
   reg _409653_409653 ; 
   reg __409653_409653;
   reg _409654_409654 ; 
   reg __409654_409654;
   reg _409655_409655 ; 
   reg __409655_409655;
   reg _409656_409656 ; 
   reg __409656_409656;
   reg _409657_409657 ; 
   reg __409657_409657;
   reg _409658_409658 ; 
   reg __409658_409658;
   reg _409659_409659 ; 
   reg __409659_409659;
   reg _409660_409660 ; 
   reg __409660_409660;
   reg _409661_409661 ; 
   reg __409661_409661;
   reg _409662_409662 ; 
   reg __409662_409662;
   reg _409663_409663 ; 
   reg __409663_409663;
   reg _409664_409664 ; 
   reg __409664_409664;
   reg _409665_409665 ; 
   reg __409665_409665;
   reg _409666_409666 ; 
   reg __409666_409666;
   reg _409667_409667 ; 
   reg __409667_409667;
   reg _409668_409668 ; 
   reg __409668_409668;
   reg _409669_409669 ; 
   reg __409669_409669;
   reg _409670_409670 ; 
   reg __409670_409670;
   reg _409671_409671 ; 
   reg __409671_409671;
   reg _409672_409672 ; 
   reg __409672_409672;
   reg _409673_409673 ; 
   reg __409673_409673;
   reg _409674_409674 ; 
   reg __409674_409674;
   reg _409675_409675 ; 
   reg __409675_409675;
   reg _409676_409676 ; 
   reg __409676_409676;
   reg _409677_409677 ; 
   reg __409677_409677;
   reg _409678_409678 ; 
   reg __409678_409678;
   reg _409679_409679 ; 
   reg __409679_409679;
   reg _409680_409680 ; 
   reg __409680_409680;
   reg _409681_409681 ; 
   reg __409681_409681;
   reg _409682_409682 ; 
   reg __409682_409682;
   reg _409683_409683 ; 
   reg __409683_409683;
   reg _409684_409684 ; 
   reg __409684_409684;
   reg _409685_409685 ; 
   reg __409685_409685;
   reg _409686_409686 ; 
   reg __409686_409686;
   reg _409687_409687 ; 
   reg __409687_409687;
   reg _409688_409688 ; 
   reg __409688_409688;
   reg _409689_409689 ; 
   reg __409689_409689;
   reg _409690_409690 ; 
   reg __409690_409690;
   reg _409691_409691 ; 
   reg __409691_409691;
   reg _409692_409692 ; 
   reg __409692_409692;
   reg _409693_409693 ; 
   reg __409693_409693;
   reg _409694_409694 ; 
   reg __409694_409694;
   reg _409695_409695 ; 
   reg __409695_409695;
   reg _409696_409696 ; 
   reg __409696_409696;
   reg _409697_409697 ; 
   reg __409697_409697;
   reg _409698_409698 ; 
   reg __409698_409698;
   reg _409699_409699 ; 
   reg __409699_409699;
   reg _409700_409700 ; 
   reg __409700_409700;
   reg _409701_409701 ; 
   reg __409701_409701;
   reg _409702_409702 ; 
   reg __409702_409702;
   reg _409703_409703 ; 
   reg __409703_409703;
   reg _409704_409704 ; 
   reg __409704_409704;
   reg _409705_409705 ; 
   reg __409705_409705;
   reg _409706_409706 ; 
   reg __409706_409706;
   reg _409707_409707 ; 
   reg __409707_409707;
   reg _409708_409708 ; 
   reg __409708_409708;
   reg _409709_409709 ; 
   reg __409709_409709;
   reg _409710_409710 ; 
   reg __409710_409710;
   reg _409711_409711 ; 
   reg __409711_409711;
   reg _409712_409712 ; 
   reg __409712_409712;
   reg _409713_409713 ; 
   reg __409713_409713;
   reg _409714_409714 ; 
   reg __409714_409714;
   reg _409715_409715 ; 
   reg __409715_409715;
   reg _409716_409716 ; 
   reg __409716_409716;
   reg _409717_409717 ; 
   reg __409717_409717;
   reg _409718_409718 ; 
   reg __409718_409718;
   reg _409719_409719 ; 
   reg __409719_409719;
   reg _409720_409720 ; 
   reg __409720_409720;
   reg _409721_409721 ; 
   reg __409721_409721;
   reg _409722_409722 ; 
   reg __409722_409722;
   reg _409723_409723 ; 
   reg __409723_409723;
   reg _409724_409724 ; 
   reg __409724_409724;
   reg _409725_409725 ; 
   reg __409725_409725;
   reg _409726_409726 ; 
   reg __409726_409726;
   reg _409727_409727 ; 
   reg __409727_409727;
   reg _409728_409728 ; 
   reg __409728_409728;
   reg _409729_409729 ; 
   reg __409729_409729;
   reg _409730_409730 ; 
   reg __409730_409730;
   reg _409731_409731 ; 
   reg __409731_409731;
   reg _409732_409732 ; 
   reg __409732_409732;
   reg _409733_409733 ; 
   reg __409733_409733;
   reg _409734_409734 ; 
   reg __409734_409734;
   reg _409735_409735 ; 
   reg __409735_409735;
   reg _409736_409736 ; 
   reg __409736_409736;
   reg _409737_409737 ; 
   reg __409737_409737;
   reg _409738_409738 ; 
   reg __409738_409738;
   reg _409739_409739 ; 
   reg __409739_409739;
   reg _409740_409740 ; 
   reg __409740_409740;
   reg _409741_409741 ; 
   reg __409741_409741;
   reg _409742_409742 ; 
   reg __409742_409742;
   reg _409743_409743 ; 
   reg __409743_409743;
   reg _409744_409744 ; 
   reg __409744_409744;
   reg _409745_409745 ; 
   reg __409745_409745;
   reg _409746_409746 ; 
   reg __409746_409746;
   reg _409747_409747 ; 
   reg __409747_409747;
   reg _409748_409748 ; 
   reg __409748_409748;
   reg _409749_409749 ; 
   reg __409749_409749;
   reg _409750_409750 ; 
   reg __409750_409750;
   reg _409751_409751 ; 
   reg __409751_409751;
   reg _409752_409752 ; 
   reg __409752_409752;
   reg _409753_409753 ; 
   reg __409753_409753;
   reg _409754_409754 ; 
   reg __409754_409754;
   reg _409755_409755 ; 
   reg __409755_409755;
   reg _409756_409756 ; 
   reg __409756_409756;
   reg _409757_409757 ; 
   reg __409757_409757;
   reg _409758_409758 ; 
   reg __409758_409758;
   reg _409759_409759 ; 
   reg __409759_409759;
   reg _409760_409760 ; 
   reg __409760_409760;
   reg _409761_409761 ; 
   reg __409761_409761;
   reg _409762_409762 ; 
   reg __409762_409762;
   reg _409763_409763 ; 
   reg __409763_409763;
   reg _409764_409764 ; 
   reg __409764_409764;
   reg _409765_409765 ; 
   reg __409765_409765;
   reg _409766_409766 ; 
   reg __409766_409766;
   reg _409767_409767 ; 
   reg __409767_409767;
   reg _409768_409768 ; 
   reg __409768_409768;
   reg _409769_409769 ; 
   reg __409769_409769;
   reg _409770_409770 ; 
   reg __409770_409770;
   reg _409771_409771 ; 
   reg __409771_409771;
   reg _409772_409772 ; 
   reg __409772_409772;
   reg _409773_409773 ; 
   reg __409773_409773;
   reg _409774_409774 ; 
   reg __409774_409774;
   reg _409775_409775 ; 
   reg __409775_409775;
   reg _409776_409776 ; 
   reg __409776_409776;
   reg _409777_409777 ; 
   reg __409777_409777;
   reg _409778_409778 ; 
   reg __409778_409778;
   reg _409779_409779 ; 
   reg __409779_409779;
   reg _409780_409780 ; 
   reg __409780_409780;
   reg _409781_409781 ; 
   reg __409781_409781;
   reg _409782_409782 ; 
   reg __409782_409782;
   reg _409783_409783 ; 
   reg __409783_409783;
   reg _409784_409784 ; 
   reg __409784_409784;
   reg _409785_409785 ; 
   reg __409785_409785;
   reg _409786_409786 ; 
   reg __409786_409786;
   reg _409787_409787 ; 
   reg __409787_409787;
   reg _409788_409788 ; 
   reg __409788_409788;
   reg _409789_409789 ; 
   reg __409789_409789;
   reg _409790_409790 ; 
   reg __409790_409790;
   reg _409791_409791 ; 
   reg __409791_409791;
   reg _409792_409792 ; 
   reg __409792_409792;
   reg _409793_409793 ; 
   reg __409793_409793;
   reg _409794_409794 ; 
   reg __409794_409794;
   reg _409795_409795 ; 
   reg __409795_409795;
   reg _409796_409796 ; 
   reg __409796_409796;
   reg _409797_409797 ; 
   reg __409797_409797;
   reg _409798_409798 ; 
   reg __409798_409798;
   reg _409799_409799 ; 
   reg __409799_409799;
   reg _409800_409800 ; 
   reg __409800_409800;
   reg _409801_409801 ; 
   reg __409801_409801;
   reg _409802_409802 ; 
   reg __409802_409802;
   reg _409803_409803 ; 
   reg __409803_409803;
   reg _409804_409804 ; 
   reg __409804_409804;
   reg _409805_409805 ; 
   reg __409805_409805;
   reg _409806_409806 ; 
   reg __409806_409806;
   reg _409807_409807 ; 
   reg __409807_409807;
   reg _409808_409808 ; 
   reg __409808_409808;
   reg _409809_409809 ; 
   reg __409809_409809;
   reg _409810_409810 ; 
   reg __409810_409810;
   reg _409811_409811 ; 
   reg __409811_409811;
   reg _409812_409812 ; 
   reg __409812_409812;
   reg _409813_409813 ; 
   reg __409813_409813;
   reg _409814_409814 ; 
   reg __409814_409814;
   reg _409815_409815 ; 
   reg __409815_409815;
   reg _409816_409816 ; 
   reg __409816_409816;
   reg _409817_409817 ; 
   reg __409817_409817;
   reg _409818_409818 ; 
   reg __409818_409818;
   reg _409819_409819 ; 
   reg __409819_409819;
   reg _409820_409820 ; 
   reg __409820_409820;
   reg _409821_409821 ; 
   reg __409821_409821;
   reg _409822_409822 ; 
   reg __409822_409822;
   reg _409823_409823 ; 
   reg __409823_409823;
   reg _409824_409824 ; 
   reg __409824_409824;
   reg _409825_409825 ; 
   reg __409825_409825;
   reg _409826_409826 ; 
   reg __409826_409826;
   reg _409827_409827 ; 
   reg __409827_409827;
   reg _409828_409828 ; 
   reg __409828_409828;
   reg _409829_409829 ; 
   reg __409829_409829;
   reg _409830_409830 ; 
   reg __409830_409830;
   reg _409831_409831 ; 
   reg __409831_409831;
   reg _409832_409832 ; 
   reg __409832_409832;
   reg _409833_409833 ; 
   reg __409833_409833;
   reg _409834_409834 ; 
   reg __409834_409834;
   reg _409835_409835 ; 
   reg __409835_409835;
   reg _409836_409836 ; 
   reg __409836_409836;
   reg _409837_409837 ; 
   reg __409837_409837;
   reg _409838_409838 ; 
   reg __409838_409838;
   reg _409839_409839 ; 
   reg __409839_409839;
   reg _409840_409840 ; 
   reg __409840_409840;
   reg _409841_409841 ; 
   reg __409841_409841;
   reg _409842_409842 ; 
   reg __409842_409842;
   reg _409843_409843 ; 
   reg __409843_409843;
   reg _409844_409844 ; 
   reg __409844_409844;
   reg _409845_409845 ; 
   reg __409845_409845;
   reg _409846_409846 ; 
   reg __409846_409846;
   reg _409847_409847 ; 
   reg __409847_409847;
   reg _409848_409848 ; 
   reg __409848_409848;
   reg _409849_409849 ; 
   reg __409849_409849;
   reg _409850_409850 ; 
   reg __409850_409850;
   reg _409851_409851 ; 
   reg __409851_409851;
   reg _409852_409852 ; 
   reg __409852_409852;
   reg _409853_409853 ; 
   reg __409853_409853;
   reg _409854_409854 ; 
   reg __409854_409854;
   reg _409855_409855 ; 
   reg __409855_409855;
   reg _409856_409856 ; 
   reg __409856_409856;
   reg _409857_409857 ; 
   reg __409857_409857;
   reg _409858_409858 ; 
   reg __409858_409858;
   reg _409859_409859 ; 
   reg __409859_409859;
   reg _409860_409860 ; 
   reg __409860_409860;
   reg _409861_409861 ; 
   reg __409861_409861;
   reg _409862_409862 ; 
   reg __409862_409862;
   reg _409863_409863 ; 
   reg __409863_409863;
   reg _409864_409864 ; 
   reg __409864_409864;
   reg _409865_409865 ; 
   reg __409865_409865;
   reg _409866_409866 ; 
   reg __409866_409866;
   reg _409867_409867 ; 
   reg __409867_409867;
   reg _409868_409868 ; 
   reg __409868_409868;
   reg _409869_409869 ; 
   reg __409869_409869;
   reg _409870_409870 ; 
   reg __409870_409870;
   reg _409871_409871 ; 
   reg __409871_409871;
   reg _409872_409872 ; 
   reg __409872_409872;
   reg _409873_409873 ; 
   reg __409873_409873;
   reg _409874_409874 ; 
   reg __409874_409874;
   reg _409875_409875 ; 
   reg __409875_409875;
   reg _409876_409876 ; 
   reg __409876_409876;
   reg _409877_409877 ; 
   reg __409877_409877;
   reg _409878_409878 ; 
   reg __409878_409878;
   reg _409879_409879 ; 
   reg __409879_409879;
   reg _409880_409880 ; 
   reg __409880_409880;
   reg _409881_409881 ; 
   reg __409881_409881;
   reg _409882_409882 ; 
   reg __409882_409882;
   reg _409883_409883 ; 
   reg __409883_409883;
   reg _409884_409884 ; 
   reg __409884_409884;
   reg _409885_409885 ; 
   reg __409885_409885;
   reg _409886_409886 ; 
   reg __409886_409886;
   reg _409887_409887 ; 
   reg __409887_409887;
   reg _409888_409888 ; 
   reg __409888_409888;
   reg _409889_409889 ; 
   reg __409889_409889;
   reg _409890_409890 ; 
   reg __409890_409890;
   reg _409891_409891 ; 
   reg __409891_409891;
   reg _409892_409892 ; 
   reg __409892_409892;
   reg _409893_409893 ; 
   reg __409893_409893;
   reg _409894_409894 ; 
   reg __409894_409894;
   reg _409895_409895 ; 
   reg __409895_409895;
   reg _409896_409896 ; 
   reg __409896_409896;
   reg _409897_409897 ; 
   reg __409897_409897;
   reg _409898_409898 ; 
   reg __409898_409898;
   reg _409899_409899 ; 
   reg __409899_409899;
   reg _409900_409900 ; 
   reg __409900_409900;
   reg _409901_409901 ; 
   reg __409901_409901;
   reg _409902_409902 ; 
   reg __409902_409902;
   reg _409903_409903 ; 
   reg __409903_409903;
   reg _409904_409904 ; 
   reg __409904_409904;
   reg _409905_409905 ; 
   reg __409905_409905;
   reg _409906_409906 ; 
   reg __409906_409906;
   reg _409907_409907 ; 
   reg __409907_409907;
   reg _409908_409908 ; 
   reg __409908_409908;
   reg _409909_409909 ; 
   reg __409909_409909;
   reg _409910_409910 ; 
   reg __409910_409910;
   reg _409911_409911 ; 
   reg __409911_409911;
   reg _409912_409912 ; 
   reg __409912_409912;
   reg _409913_409913 ; 
   reg __409913_409913;
   reg _409914_409914 ; 
   reg __409914_409914;
   reg _409915_409915 ; 
   reg __409915_409915;
   reg _409916_409916 ; 
   reg __409916_409916;
   reg _409917_409917 ; 
   reg __409917_409917;
   reg _409918_409918 ; 
   reg __409918_409918;
   reg _409919_409919 ; 
   reg __409919_409919;
   reg _409920_409920 ; 
   reg __409920_409920;
   reg _409921_409921 ; 
   reg __409921_409921;
   reg _409922_409922 ; 
   reg __409922_409922;
   reg _409923_409923 ; 
   reg __409923_409923;
   reg _409924_409924 ; 
   reg __409924_409924;
   reg _409925_409925 ; 
   reg __409925_409925;
   reg _409926_409926 ; 
   reg __409926_409926;
   reg _409927_409927 ; 
   reg __409927_409927;
   reg _409928_409928 ; 
   reg __409928_409928;
   reg _409929_409929 ; 
   reg __409929_409929;
   reg _409930_409930 ; 
   reg __409930_409930;
   reg _409931_409931 ; 
   reg __409931_409931;
   reg _409932_409932 ; 
   reg __409932_409932;
   reg _409933_409933 ; 
   reg __409933_409933;
   reg _409934_409934 ; 
   reg __409934_409934;
   reg _409935_409935 ; 
   reg __409935_409935;
   reg _409936_409936 ; 
   reg __409936_409936;
   reg _409937_409937 ; 
   reg __409937_409937;
   reg _409938_409938 ; 
   reg __409938_409938;
   reg _409939_409939 ; 
   reg __409939_409939;
   reg _409940_409940 ; 
   reg __409940_409940;
   reg _409941_409941 ; 
   reg __409941_409941;
   reg _409942_409942 ; 
   reg __409942_409942;
   reg _409943_409943 ; 
   reg __409943_409943;
   reg _409944_409944 ; 
   reg __409944_409944;
   reg _409945_409945 ; 
   reg __409945_409945;
   reg _409946_409946 ; 
   reg __409946_409946;
   reg _409947_409947 ; 
   reg __409947_409947;
   reg _409948_409948 ; 
   reg __409948_409948;
   reg _409949_409949 ; 
   reg __409949_409949;
   reg _409950_409950 ; 
   reg __409950_409950;
   reg _409951_409951 ; 
   reg __409951_409951;
   reg _409952_409952 ; 
   reg __409952_409952;
   reg _409953_409953 ; 
   reg __409953_409953;
   reg _409954_409954 ; 
   reg __409954_409954;
   reg _409955_409955 ; 
   reg __409955_409955;
   reg _409956_409956 ; 
   reg __409956_409956;
   reg _409957_409957 ; 
   reg __409957_409957;
   reg _409958_409958 ; 
   reg __409958_409958;
   reg _409959_409959 ; 
   reg __409959_409959;
   reg _409960_409960 ; 
   reg __409960_409960;
   reg _409961_409961 ; 
   reg __409961_409961;
   reg _409962_409962 ; 
   reg __409962_409962;
   reg _409963_409963 ; 
   reg __409963_409963;
   reg _409964_409964 ; 
   reg __409964_409964;
   reg _409965_409965 ; 
   reg __409965_409965;
   reg _409966_409966 ; 
   reg __409966_409966;
   reg _409967_409967 ; 
   reg __409967_409967;
   reg _409968_409968 ; 
   reg __409968_409968;
   reg _409969_409969 ; 
   reg __409969_409969;
   reg _409970_409970 ; 
   reg __409970_409970;
   reg _409971_409971 ; 
   reg __409971_409971;
   reg _409972_409972 ; 
   reg __409972_409972;
   reg _409973_409973 ; 
   reg __409973_409973;
   reg _409974_409974 ; 
   reg __409974_409974;
   reg _409975_409975 ; 
   reg __409975_409975;
   reg _409976_409976 ; 
   reg __409976_409976;
   reg _409977_409977 ; 
   reg __409977_409977;
   reg _409978_409978 ; 
   reg __409978_409978;
   reg _409979_409979 ; 
   reg __409979_409979;
   reg _409980_409980 ; 
   reg __409980_409980;
   reg _409981_409981 ; 
   reg __409981_409981;
   reg _409982_409982 ; 
   reg __409982_409982;
   reg _409983_409983 ; 
   reg __409983_409983;
   reg _409984_409984 ; 
   reg __409984_409984;
   reg _409985_409985 ; 
   reg __409985_409985;
   reg _409986_409986 ; 
   reg __409986_409986;
   reg _409987_409987 ; 
   reg __409987_409987;
   reg _409988_409988 ; 
   reg __409988_409988;
   reg _409989_409989 ; 
   reg __409989_409989;
   reg _409990_409990 ; 
   reg __409990_409990;
   reg _409991_409991 ; 
   reg __409991_409991;
   reg _409992_409992 ; 
   reg __409992_409992;
   reg _409993_409993 ; 
   reg __409993_409993;
   reg _409994_409994 ; 
   reg __409994_409994;
   reg _409995_409995 ; 
   reg __409995_409995;
   reg _409996_409996 ; 
   reg __409996_409996;
   reg _409997_409997 ; 
   reg __409997_409997;
   reg _409998_409998 ; 
   reg __409998_409998;
   reg _409999_409999 ; 
   reg __409999_409999;
   reg _410000_410000 ; 
   reg __410000_410000;
   reg _410001_410001 ; 
   reg __410001_410001;
   reg _410002_410002 ; 
   reg __410002_410002;
   reg _410003_410003 ; 
   reg __410003_410003;
   reg _410004_410004 ; 
   reg __410004_410004;
   reg _410005_410005 ; 
   reg __410005_410005;
   reg _410006_410006 ; 
   reg __410006_410006;
   reg _410007_410007 ; 
   reg __410007_410007;
   reg _410008_410008 ; 
   reg __410008_410008;
   reg _410009_410009 ; 
   reg __410009_410009;
   reg _410010_410010 ; 
   reg __410010_410010;
   reg _410011_410011 ; 
   reg __410011_410011;
   reg _410012_410012 ; 
   reg __410012_410012;
   reg _410013_410013 ; 
   reg __410013_410013;
   reg _410014_410014 ; 
   reg __410014_410014;
   reg _410015_410015 ; 
   reg __410015_410015;
   reg _410016_410016 ; 
   reg __410016_410016;
   reg _410017_410017 ; 
   reg __410017_410017;
   reg _410018_410018 ; 
   reg __410018_410018;
   reg _410019_410019 ; 
   reg __410019_410019;
   reg _410020_410020 ; 
   reg __410020_410020;
   reg _410021_410021 ; 
   reg __410021_410021;
   reg _410022_410022 ; 
   reg __410022_410022;
   reg _410023_410023 ; 
   reg __410023_410023;
   reg _410024_410024 ; 
   reg __410024_410024;
   reg _410025_410025 ; 
   reg __410025_410025;
   reg _410026_410026 ; 
   reg __410026_410026;
   reg _410027_410027 ; 
   reg __410027_410027;
   reg _410028_410028 ; 
   reg __410028_410028;
   reg _410029_410029 ; 
   reg __410029_410029;
   reg _410030_410030 ; 
   reg __410030_410030;
   reg _410031_410031 ; 
   reg __410031_410031;
   reg _410032_410032 ; 
   reg __410032_410032;
   reg _410033_410033 ; 
   reg __410033_410033;
   reg _410034_410034 ; 
   reg __410034_410034;
   reg _410035_410035 ; 
   reg __410035_410035;
   reg _410036_410036 ; 
   reg __410036_410036;
   reg _410037_410037 ; 
   reg __410037_410037;
   reg _410038_410038 ; 
   reg __410038_410038;
   reg _410039_410039 ; 
   reg __410039_410039;
   reg _410040_410040 ; 
   reg __410040_410040;
   reg _410041_410041 ; 
   reg __410041_410041;
   reg _410042_410042 ; 
   reg __410042_410042;
   reg _410043_410043 ; 
   reg __410043_410043;
   reg _410044_410044 ; 
   reg __410044_410044;
   reg _410045_410045 ; 
   reg __410045_410045;
   reg _410046_410046 ; 
   reg __410046_410046;
   reg _410047_410047 ; 
   reg __410047_410047;
   reg _410048_410048 ; 
   reg __410048_410048;
   reg _410049_410049 ; 
   reg __410049_410049;
   reg _410050_410050 ; 
   reg __410050_410050;
   reg _410051_410051 ; 
   reg __410051_410051;
   reg _410052_410052 ; 
   reg __410052_410052;
   reg _410053_410053 ; 
   reg __410053_410053;
   reg _410054_410054 ; 
   reg __410054_410054;
   reg _410055_410055 ; 
   reg __410055_410055;
   reg _410056_410056 ; 
   reg __410056_410056;
   reg _410057_410057 ; 
   reg __410057_410057;
   reg _410058_410058 ; 
   reg __410058_410058;
   reg _410059_410059 ; 
   reg __410059_410059;
   reg _410060_410060 ; 
   reg __410060_410060;
   reg _410061_410061 ; 
   reg __410061_410061;
   reg _410062_410062 ; 
   reg __410062_410062;
   reg _410063_410063 ; 
   reg __410063_410063;
   reg _410064_410064 ; 
   reg __410064_410064;
   reg _410065_410065 ; 
   reg __410065_410065;
   reg _410066_410066 ; 
   reg __410066_410066;
   reg _410067_410067 ; 
   reg __410067_410067;
   reg _410068_410068 ; 
   reg __410068_410068;
   reg _410069_410069 ; 
   reg __410069_410069;
   reg _410070_410070 ; 
   reg __410070_410070;
   reg _410071_410071 ; 
   reg __410071_410071;
   reg _410072_410072 ; 
   reg __410072_410072;
   reg _410073_410073 ; 
   reg __410073_410073;
   reg _410074_410074 ; 
   reg __410074_410074;
   reg _410075_410075 ; 
   reg __410075_410075;
   reg _410076_410076 ; 
   reg __410076_410076;
   reg _410077_410077 ; 
   reg __410077_410077;
   reg _410078_410078 ; 
   reg __410078_410078;
   reg _410079_410079 ; 
   reg __410079_410079;
   reg _410080_410080 ; 
   reg __410080_410080;
   reg _410081_410081 ; 
   reg __410081_410081;
   reg _410082_410082 ; 
   reg __410082_410082;
   reg _410083_410083 ; 
   reg __410083_410083;
   reg _410084_410084 ; 
   reg __410084_410084;
   reg _410085_410085 ; 
   reg __410085_410085;
   reg _410086_410086 ; 
   reg __410086_410086;
   reg _410087_410087 ; 
   reg __410087_410087;
   reg _410088_410088 ; 
   reg __410088_410088;
   reg _410089_410089 ; 
   reg __410089_410089;
   reg _410090_410090 ; 
   reg __410090_410090;
   reg _410091_410091 ; 
   reg __410091_410091;
   reg _410092_410092 ; 
   reg __410092_410092;
   reg _410093_410093 ; 
   reg __410093_410093;
   reg _410094_410094 ; 
   reg __410094_410094;
   reg _410095_410095 ; 
   reg __410095_410095;
   reg _410096_410096 ; 
   reg __410096_410096;
   reg _410097_410097 ; 
   reg __410097_410097;
   reg _410098_410098 ; 
   reg __410098_410098;
   reg _410099_410099 ; 
   reg __410099_410099;
   reg _410100_410100 ; 
   reg __410100_410100;
   reg _410101_410101 ; 
   reg __410101_410101;
   reg _410102_410102 ; 
   reg __410102_410102;
   reg _410103_410103 ; 
   reg __410103_410103;
   reg _410104_410104 ; 
   reg __410104_410104;
   reg _410105_410105 ; 
   reg __410105_410105;
   reg _410106_410106 ; 
   reg __410106_410106;
   reg _410107_410107 ; 
   reg __410107_410107;
   reg _410108_410108 ; 
   reg __410108_410108;
   reg _410109_410109 ; 
   reg __410109_410109;
   reg _410110_410110 ; 
   reg __410110_410110;
   reg _410111_410111 ; 
   reg __410111_410111;
   reg _410112_410112 ; 
   reg __410112_410112;
   reg _410113_410113 ; 
   reg __410113_410113;
   reg _410114_410114 ; 
   reg __410114_410114;
   reg _410115_410115 ; 
   reg __410115_410115;
   reg _410116_410116 ; 
   reg __410116_410116;
   reg _410117_410117 ; 
   reg __410117_410117;
   reg _410118_410118 ; 
   reg __410118_410118;
   reg _410119_410119 ; 
   reg __410119_410119;
   reg _410120_410120 ; 
   reg __410120_410120;
   reg _410121_410121 ; 
   reg __410121_410121;
   reg _410122_410122 ; 
   reg __410122_410122;
   reg _410123_410123 ; 
   reg __410123_410123;
   reg _410124_410124 ; 
   reg __410124_410124;
   reg _410125_410125 ; 
   reg __410125_410125;
   reg _410126_410126 ; 
   reg __410126_410126;
   reg _410127_410127 ; 
   reg __410127_410127;
   reg _410128_410128 ; 
   reg __410128_410128;
   reg _410129_410129 ; 
   reg __410129_410129;
   reg _410130_410130 ; 
   reg __410130_410130;
   reg _410131_410131 ; 
   reg __410131_410131;
   reg _410132_410132 ; 
   reg __410132_410132;
   reg _410133_410133 ; 
   reg __410133_410133;
   reg _410134_410134 ; 
   reg __410134_410134;
   reg _410135_410135 ; 
   reg __410135_410135;
   reg _410136_410136 ; 
   reg __410136_410136;
   reg _410137_410137 ; 
   reg __410137_410137;
   reg _410138_410138 ; 
   reg __410138_410138;
   reg _410139_410139 ; 
   reg __410139_410139;
   reg _410140_410140 ; 
   reg __410140_410140;
   reg _410141_410141 ; 
   reg __410141_410141;
   reg _410142_410142 ; 
   reg __410142_410142;
   reg _410143_410143 ; 
   reg __410143_410143;
   reg _410144_410144 ; 
   reg __410144_410144;
   reg _410145_410145 ; 
   reg __410145_410145;
   reg _410146_410146 ; 
   reg __410146_410146;
   reg _410147_410147 ; 
   reg __410147_410147;
   reg _410148_410148 ; 
   reg __410148_410148;
   reg _410149_410149 ; 
   reg __410149_410149;
   reg _410150_410150 ; 
   reg __410150_410150;
   reg _410151_410151 ; 
   reg __410151_410151;
   reg _410152_410152 ; 
   reg __410152_410152;
   reg _410153_410153 ; 
   reg __410153_410153;
   reg _410154_410154 ; 
   reg __410154_410154;
   reg _410155_410155 ; 
   reg __410155_410155;
   reg _410156_410156 ; 
   reg __410156_410156;
   reg _410157_410157 ; 
   reg __410157_410157;
   reg _410158_410158 ; 
   reg __410158_410158;
   reg _410159_410159 ; 
   reg __410159_410159;
   reg _410160_410160 ; 
   reg __410160_410160;
   reg _410161_410161 ; 
   reg __410161_410161;
   reg _410162_410162 ; 
   reg __410162_410162;
   reg _410163_410163 ; 
   reg __410163_410163;
   reg _410164_410164 ; 
   reg __410164_410164;
   reg _410165_410165 ; 
   reg __410165_410165;
   reg _410166_410166 ; 
   reg __410166_410166;
   reg _410167_410167 ; 
   reg __410167_410167;
   reg _410168_410168 ; 
   reg __410168_410168;
   reg _410169_410169 ; 
   reg __410169_410169;
   reg _410170_410170 ; 
   reg __410170_410170;
   reg _410171_410171 ; 
   reg __410171_410171;
   reg _410172_410172 ; 
   reg __410172_410172;
   reg _410173_410173 ; 
   reg __410173_410173;
   reg _410174_410174 ; 
   reg __410174_410174;
   reg _410175_410175 ; 
   reg __410175_410175;
   reg _410176_410176 ; 
   reg __410176_410176;
   reg _410177_410177 ; 
   reg __410177_410177;
   reg _410178_410178 ; 
   reg __410178_410178;
   reg _410179_410179 ; 
   reg __410179_410179;
   reg _410180_410180 ; 
   reg __410180_410180;
   reg _410181_410181 ; 
   reg __410181_410181;
   reg _410182_410182 ; 
   reg __410182_410182;
   reg _410183_410183 ; 
   reg __410183_410183;
   reg _410184_410184 ; 
   reg __410184_410184;
   reg _410185_410185 ; 
   reg __410185_410185;
   reg _410186_410186 ; 
   reg __410186_410186;
   reg _410187_410187 ; 
   reg __410187_410187;
   reg _410188_410188 ; 
   reg __410188_410188;
   reg _410189_410189 ; 
   reg __410189_410189;
   reg _410190_410190 ; 
   reg __410190_410190;
   reg _410191_410191 ; 
   reg __410191_410191;
   reg _410192_410192 ; 
   reg __410192_410192;
   reg _410193_410193 ; 
   reg __410193_410193;
   reg _410194_410194 ; 
   reg __410194_410194;
   reg _410195_410195 ; 
   reg __410195_410195;
   reg _410196_410196 ; 
   reg __410196_410196;
   reg _410197_410197 ; 
   reg __410197_410197;
   reg _410198_410198 ; 
   reg __410198_410198;
   reg _410199_410199 ; 
   reg __410199_410199;
   reg _410200_410200 ; 
   reg __410200_410200;
   reg _410201_410201 ; 
   reg __410201_410201;
   reg _410202_410202 ; 
   reg __410202_410202;
   reg _410203_410203 ; 
   reg __410203_410203;
   reg _410204_410204 ; 
   reg __410204_410204;
   reg _410205_410205 ; 
   reg __410205_410205;
   reg _410206_410206 ; 
   reg __410206_410206;
   reg _410207_410207 ; 
   reg __410207_410207;
   reg _410208_410208 ; 
   reg __410208_410208;
   reg _410209_410209 ; 
   reg __410209_410209;
   reg _410210_410210 ; 
   reg __410210_410210;
   reg _410211_410211 ; 
   reg __410211_410211;
   reg _410212_410212 ; 
   reg __410212_410212;
   reg _410213_410213 ; 
   reg __410213_410213;
   reg _410214_410214 ; 
   reg __410214_410214;
   reg _410215_410215 ; 
   reg __410215_410215;
   reg _410216_410216 ; 
   reg __410216_410216;
   reg _410217_410217 ; 
   reg __410217_410217;
   reg _410218_410218 ; 
   reg __410218_410218;
   reg _410219_410219 ; 
   reg __410219_410219;
   reg _410220_410220 ; 
   reg __410220_410220;
   reg _410221_410221 ; 
   reg __410221_410221;
   reg _410222_410222 ; 
   reg __410222_410222;
   reg _410223_410223 ; 
   reg __410223_410223;
   reg _410224_410224 ; 
   reg __410224_410224;
   reg _410225_410225 ; 
   reg __410225_410225;
   reg _410226_410226 ; 
   reg __410226_410226;
   reg _410227_410227 ; 
   reg __410227_410227;
   reg _410228_410228 ; 
   reg __410228_410228;
   reg _410229_410229 ; 
   reg __410229_410229;
   reg _410230_410230 ; 
   reg __410230_410230;
   reg _410231_410231 ; 
   reg __410231_410231;
   reg _410232_410232 ; 
   reg __410232_410232;
   reg _410233_410233 ; 
   reg __410233_410233;
   reg _410234_410234 ; 
   reg __410234_410234;
   reg _410235_410235 ; 
   reg __410235_410235;
   reg _410236_410236 ; 
   reg __410236_410236;
   reg _410237_410237 ; 
   reg __410237_410237;
   reg _410238_410238 ; 
   reg __410238_410238;
   reg _410239_410239 ; 
   reg __410239_410239;
   reg _410240_410240 ; 
   reg __410240_410240;
   reg _410241_410241 ; 
   reg __410241_410241;
   reg _410242_410242 ; 
   reg __410242_410242;
   reg _410243_410243 ; 
   reg __410243_410243;
   reg _410244_410244 ; 
   reg __410244_410244;
   reg _410245_410245 ; 
   reg __410245_410245;
   reg _410246_410246 ; 
   reg __410246_410246;
   reg _410247_410247 ; 
   reg __410247_410247;
   reg _410248_410248 ; 
   reg __410248_410248;
   reg _410249_410249 ; 
   reg __410249_410249;
   reg _410250_410250 ; 
   reg __410250_410250;
   reg _410251_410251 ; 
   reg __410251_410251;
   reg _410252_410252 ; 
   reg __410252_410252;
   reg _410253_410253 ; 
   reg __410253_410253;
   reg _410254_410254 ; 
   reg __410254_410254;
   reg _410255_410255 ; 
   reg __410255_410255;
   reg _410256_410256 ; 
   reg __410256_410256;
   reg _410257_410257 ; 
   reg __410257_410257;
   reg _410258_410258 ; 
   reg __410258_410258;
   reg _410259_410259 ; 
   reg __410259_410259;
   reg _410260_410260 ; 
   reg __410260_410260;
   reg _410261_410261 ; 
   reg __410261_410261;
   reg _410262_410262 ; 
   reg __410262_410262;
   reg _410263_410263 ; 
   reg __410263_410263;
   reg _410264_410264 ; 
   reg __410264_410264;
   reg _410265_410265 ; 
   reg __410265_410265;
   reg _410266_410266 ; 
   reg __410266_410266;
   reg _410267_410267 ; 
   reg __410267_410267;
   reg _410268_410268 ; 
   reg __410268_410268;
   reg _410269_410269 ; 
   reg __410269_410269;
   reg _410270_410270 ; 
   reg __410270_410270;
   reg _410271_410271 ; 
   reg __410271_410271;
   reg _410272_410272 ; 
   reg __410272_410272;
   reg _410273_410273 ; 
   reg __410273_410273;
   reg _410274_410274 ; 
   reg __410274_410274;
   reg _410275_410275 ; 
   reg __410275_410275;
   reg _410276_410276 ; 
   reg __410276_410276;
   reg _410277_410277 ; 
   reg __410277_410277;
   reg _410278_410278 ; 
   reg __410278_410278;
   reg _410279_410279 ; 
   reg __410279_410279;
   reg _410280_410280 ; 
   reg __410280_410280;
   reg _410281_410281 ; 
   reg __410281_410281;
   reg _410282_410282 ; 
   reg __410282_410282;
   reg _410283_410283 ; 
   reg __410283_410283;
   reg _410284_410284 ; 
   reg __410284_410284;
   reg _410285_410285 ; 
   reg __410285_410285;
   reg _410286_410286 ; 
   reg __410286_410286;
   reg _410287_410287 ; 
   reg __410287_410287;
   reg _410288_410288 ; 
   reg __410288_410288;
   reg _410289_410289 ; 
   reg __410289_410289;
   reg _410290_410290 ; 
   reg __410290_410290;
   reg _410291_410291 ; 
   reg __410291_410291;
   reg _410292_410292 ; 
   reg __410292_410292;
   reg _410293_410293 ; 
   reg __410293_410293;
   reg _410294_410294 ; 
   reg __410294_410294;
   reg _410295_410295 ; 
   reg __410295_410295;
   reg _410296_410296 ; 
   reg __410296_410296;
   reg _410297_410297 ; 
   reg __410297_410297;
   reg _410298_410298 ; 
   reg __410298_410298;
   reg _410299_410299 ; 
   reg __410299_410299;
   reg _410300_410300 ; 
   reg __410300_410300;
   reg _410301_410301 ; 
   reg __410301_410301;
   reg _410302_410302 ; 
   reg __410302_410302;
   reg _410303_410303 ; 
   reg __410303_410303;
   reg _410304_410304 ; 
   reg __410304_410304;
   reg _410305_410305 ; 
   reg __410305_410305;
   reg _410306_410306 ; 
   reg __410306_410306;
   reg _410307_410307 ; 
   reg __410307_410307;
   reg _410308_410308 ; 
   reg __410308_410308;
   reg _410309_410309 ; 
   reg __410309_410309;
   reg _410310_410310 ; 
   reg __410310_410310;
   reg _410311_410311 ; 
   reg __410311_410311;
   reg _410312_410312 ; 
   reg __410312_410312;
   reg _410313_410313 ; 
   reg __410313_410313;
   reg _410314_410314 ; 
   reg __410314_410314;
   reg _410315_410315 ; 
   reg __410315_410315;
   reg _410316_410316 ; 
   reg __410316_410316;
   reg _410317_410317 ; 
   reg __410317_410317;
   reg _410318_410318 ; 
   reg __410318_410318;
   reg _410319_410319 ; 
   reg __410319_410319;
   reg _410320_410320 ; 
   reg __410320_410320;
   reg _410321_410321 ; 
   reg __410321_410321;
   reg _410322_410322 ; 
   reg __410322_410322;
   reg _410323_410323 ; 
   reg __410323_410323;
   reg _410324_410324 ; 
   reg __410324_410324;
   reg _410325_410325 ; 
   reg __410325_410325;
   reg _410326_410326 ; 
   reg __410326_410326;
   reg _410327_410327 ; 
   reg __410327_410327;
   reg _410328_410328 ; 
   reg __410328_410328;
   reg _410329_410329 ; 
   reg __410329_410329;
   reg _410330_410330 ; 
   reg __410330_410330;
   reg _410331_410331 ; 
   reg __410331_410331;
   reg _410332_410332 ; 
   reg __410332_410332;
   reg _410333_410333 ; 
   reg __410333_410333;
   reg _410334_410334 ; 
   reg __410334_410334;
   reg _410335_410335 ; 
   reg __410335_410335;
   reg _410336_410336 ; 
   reg __410336_410336;
   reg _410337_410337 ; 
   reg __410337_410337;
   reg _410338_410338 ; 
   reg __410338_410338;
   reg _410339_410339 ; 
   reg __410339_410339;
   reg _410340_410340 ; 
   reg __410340_410340;
   reg _410341_410341 ; 
   reg __410341_410341;
   reg _410342_410342 ; 
   reg __410342_410342;
   reg _410343_410343 ; 
   reg __410343_410343;
   reg _410344_410344 ; 
   reg __410344_410344;
   reg _410345_410345 ; 
   reg __410345_410345;
   reg _410346_410346 ; 
   reg __410346_410346;
   reg _410347_410347 ; 
   reg __410347_410347;
   reg _410348_410348 ; 
   reg __410348_410348;
   reg _410349_410349 ; 
   reg __410349_410349;
   reg _410350_410350 ; 
   reg __410350_410350;
   reg _410351_410351 ; 
   reg __410351_410351;
   reg _410352_410352 ; 
   reg __410352_410352;
   reg _410353_410353 ; 
   reg __410353_410353;
   reg _410354_410354 ; 
   reg __410354_410354;
   reg _410355_410355 ; 
   reg __410355_410355;
   reg _410356_410356 ; 
   reg __410356_410356;
   reg _410357_410357 ; 
   reg __410357_410357;
   reg _410358_410358 ; 
   reg __410358_410358;
   reg _410359_410359 ; 
   reg __410359_410359;
   reg _410360_410360 ; 
   reg __410360_410360;
   reg _410361_410361 ; 
   reg __410361_410361;
   reg _410362_410362 ; 
   reg __410362_410362;
   reg _410363_410363 ; 
   reg __410363_410363;
   reg _410364_410364 ; 
   reg __410364_410364;
   reg _410365_410365 ; 
   reg __410365_410365;
   reg _410366_410366 ; 
   reg __410366_410366;
   reg _410367_410367 ; 
   reg __410367_410367;
   reg _410368_410368 ; 
   reg __410368_410368;
   reg _410369_410369 ; 
   reg __410369_410369;
   reg _410370_410370 ; 
   reg __410370_410370;
   reg _410371_410371 ; 
   reg __410371_410371;
   reg _410372_410372 ; 
   reg __410372_410372;
   reg _410373_410373 ; 
   reg __410373_410373;
   reg _410374_410374 ; 
   reg __410374_410374;
   reg _410375_410375 ; 
   reg __410375_410375;
   reg _410376_410376 ; 
   reg __410376_410376;
   reg _410377_410377 ; 
   reg __410377_410377;
   reg _410378_410378 ; 
   reg __410378_410378;
   reg _410379_410379 ; 
   reg __410379_410379;
   reg _410380_410380 ; 
   reg __410380_410380;
   reg _410381_410381 ; 
   reg __410381_410381;
   reg _410382_410382 ; 
   reg __410382_410382;
   reg _410383_410383 ; 
   reg __410383_410383;
   reg _410384_410384 ; 
   reg __410384_410384;
   reg _410385_410385 ; 
   reg __410385_410385;
   reg _410386_410386 ; 
   reg __410386_410386;
   reg _410387_410387 ; 
   reg __410387_410387;
   reg _410388_410388 ; 
   reg __410388_410388;
   reg _410389_410389 ; 
   reg __410389_410389;
   reg _410390_410390 ; 
   reg __410390_410390;
   reg _410391_410391 ; 
   reg __410391_410391;
   reg _410392_410392 ; 
   reg __410392_410392;
   reg _410393_410393 ; 
   reg __410393_410393;
   reg _410394_410394 ; 
   reg __410394_410394;
   reg _410395_410395 ; 
   reg __410395_410395;
   reg _410396_410396 ; 
   reg __410396_410396;
   reg _410397_410397 ; 
   reg __410397_410397;
   reg _410398_410398 ; 
   reg __410398_410398;
   reg _410399_410399 ; 
   reg __410399_410399;
   reg _410400_410400 ; 
   reg __410400_410400;
   reg _410401_410401 ; 
   reg __410401_410401;
   reg _410402_410402 ; 
   reg __410402_410402;
   reg _410403_410403 ; 
   reg __410403_410403;
   reg _410404_410404 ; 
   reg __410404_410404;
   reg _410405_410405 ; 
   reg __410405_410405;
   reg _410406_410406 ; 
   reg __410406_410406;
   reg _410407_410407 ; 
   reg __410407_410407;
   reg _410408_410408 ; 
   reg __410408_410408;
   reg _410409_410409 ; 
   reg __410409_410409;
   reg _410410_410410 ; 
   reg __410410_410410;
   reg _410411_410411 ; 
   reg __410411_410411;
   reg _410412_410412 ; 
   reg __410412_410412;
   reg _410413_410413 ; 
   reg __410413_410413;
   reg _410414_410414 ; 
   reg __410414_410414;
   reg _410415_410415 ; 
   reg __410415_410415;
   reg _410416_410416 ; 
   reg __410416_410416;
   reg _410417_410417 ; 
   reg __410417_410417;
   reg _410418_410418 ; 
   reg __410418_410418;
   reg _410419_410419 ; 
   reg __410419_410419;
   reg _410420_410420 ; 
   reg __410420_410420;
   reg _410421_410421 ; 
   reg __410421_410421;
   reg _410422_410422 ; 
   reg __410422_410422;
   reg _410423_410423 ; 
   reg __410423_410423;
   reg _410424_410424 ; 
   reg __410424_410424;
   reg _410425_410425 ; 
   reg __410425_410425;
   reg _410426_410426 ; 
   reg __410426_410426;
   reg _410427_410427 ; 
   reg __410427_410427;
   reg _410428_410428 ; 
   reg __410428_410428;
   reg _410429_410429 ; 
   reg __410429_410429;
   reg _410430_410430 ; 
   reg __410430_410430;
   reg _410431_410431 ; 
   reg __410431_410431;
   reg _410432_410432 ; 
   reg __410432_410432;
   reg _410433_410433 ; 
   reg __410433_410433;
   reg _410434_410434 ; 
   reg __410434_410434;
   reg _410435_410435 ; 
   reg __410435_410435;
   reg _410436_410436 ; 
   reg __410436_410436;
   reg _410437_410437 ; 
   reg __410437_410437;
   reg _410438_410438 ; 
   reg __410438_410438;
   reg _410439_410439 ; 
   reg __410439_410439;
   reg _410440_410440 ; 
   reg __410440_410440;
   reg _410441_410441 ; 
   reg __410441_410441;
   reg _410442_410442 ; 
   reg __410442_410442;
   reg _410443_410443 ; 
   reg __410443_410443;
   reg _410444_410444 ; 
   reg __410444_410444;
   reg _410445_410445 ; 
   reg __410445_410445;
   reg _410446_410446 ; 
   reg __410446_410446;
   reg _410447_410447 ; 
   reg __410447_410447;
   reg _410448_410448 ; 
   reg __410448_410448;
   reg _410449_410449 ; 
   reg __410449_410449;
   reg _410450_410450 ; 
   reg __410450_410450;
   reg _410451_410451 ; 
   reg __410451_410451;
   reg _410452_410452 ; 
   reg __410452_410452;
   reg _410453_410453 ; 
   reg __410453_410453;
   reg _410454_410454 ; 
   reg __410454_410454;
   reg _410455_410455 ; 
   reg __410455_410455;
   reg _410456_410456 ; 
   reg __410456_410456;
   reg _410457_410457 ; 
   reg __410457_410457;
   reg _410458_410458 ; 
   reg __410458_410458;
   reg _410459_410459 ; 
   reg __410459_410459;
   reg _410460_410460 ; 
   reg __410460_410460;
   reg _410461_410461 ; 
   reg __410461_410461;
   reg _410462_410462 ; 
   reg __410462_410462;
   reg _410463_410463 ; 
   reg __410463_410463;
   reg _410464_410464 ; 
   reg __410464_410464;
   reg _410465_410465 ; 
   reg __410465_410465;
   reg _410466_410466 ; 
   reg __410466_410466;
   reg _410467_410467 ; 
   reg __410467_410467;
   reg _410468_410468 ; 
   reg __410468_410468;
   reg _410469_410469 ; 
   reg __410469_410469;
   reg _410470_410470 ; 
   reg __410470_410470;
   reg _410471_410471 ; 
   reg __410471_410471;
   reg _410472_410472 ; 
   reg __410472_410472;
   reg _410473_410473 ; 
   reg __410473_410473;
   reg _410474_410474 ; 
   reg __410474_410474;
   reg _410475_410475 ; 
   reg __410475_410475;
   reg _410476_410476 ; 
   reg __410476_410476;
   reg _410477_410477 ; 
   reg __410477_410477;
   reg _410478_410478 ; 
   reg __410478_410478;
   reg _410479_410479 ; 
   reg __410479_410479;
   reg _410480_410480 ; 
   reg __410480_410480;
   reg _410481_410481 ; 
   reg __410481_410481;
   reg _410482_410482 ; 
   reg __410482_410482;
   reg _410483_410483 ; 
   reg __410483_410483;
   reg _410484_410484 ; 
   reg __410484_410484;
   reg _410485_410485 ; 
   reg __410485_410485;
   reg _410486_410486 ; 
   reg __410486_410486;
   reg _410487_410487 ; 
   reg __410487_410487;
   reg _410488_410488 ; 
   reg __410488_410488;
   reg _410489_410489 ; 
   reg __410489_410489;
   reg _410490_410490 ; 
   reg __410490_410490;
   reg _410491_410491 ; 
   reg __410491_410491;
   reg _410492_410492 ; 
   reg __410492_410492;
   reg _410493_410493 ; 
   reg __410493_410493;
   reg _410494_410494 ; 
   reg __410494_410494;
   reg _410495_410495 ; 
   reg __410495_410495;
   reg _410496_410496 ; 
   reg __410496_410496;
   reg _410497_410497 ; 
   reg __410497_410497;
   reg _410498_410498 ; 
   reg __410498_410498;
   reg _410499_410499 ; 
   reg __410499_410499;
   reg _410500_410500 ; 
   reg __410500_410500;
   reg _410501_410501 ; 
   reg __410501_410501;
   reg _410502_410502 ; 
   reg __410502_410502;
   reg _410503_410503 ; 
   reg __410503_410503;
   reg _410504_410504 ; 
   reg __410504_410504;
   reg _410505_410505 ; 
   reg __410505_410505;
   reg _410506_410506 ; 
   reg __410506_410506;
   reg _410507_410507 ; 
   reg __410507_410507;
   reg _410508_410508 ; 
   reg __410508_410508;
   reg _410509_410509 ; 
   reg __410509_410509;
   reg _410510_410510 ; 
   reg __410510_410510;
   reg _410511_410511 ; 
   reg __410511_410511;
   reg _410512_410512 ; 
   reg __410512_410512;
   reg _410513_410513 ; 
   reg __410513_410513;
   reg _410514_410514 ; 
   reg __410514_410514;
   reg _410515_410515 ; 
   reg __410515_410515;
   reg _410516_410516 ; 
   reg __410516_410516;
   reg _410517_410517 ; 
   reg __410517_410517;
   reg _410518_410518 ; 
   reg __410518_410518;
   reg _410519_410519 ; 
   reg __410519_410519;
   reg _410520_410520 ; 
   reg __410520_410520;
   reg _410521_410521 ; 
   reg __410521_410521;
   reg _410522_410522 ; 
   reg __410522_410522;
   reg _410523_410523 ; 
   reg __410523_410523;
   reg _410524_410524 ; 
   reg __410524_410524;
   reg _410525_410525 ; 
   reg __410525_410525;
   reg _410526_410526 ; 
   reg __410526_410526;
   reg _410527_410527 ; 
   reg __410527_410527;
   reg _410528_410528 ; 
   reg __410528_410528;
   reg _410529_410529 ; 
   reg __410529_410529;
   reg _410530_410530 ; 
   reg __410530_410530;
   reg _410531_410531 ; 
   reg __410531_410531;
   reg _410532_410532 ; 
   reg __410532_410532;
   reg _410533_410533 ; 
   reg __410533_410533;
   reg _410534_410534 ; 
   reg __410534_410534;
   reg _410535_410535 ; 
   reg __410535_410535;
   reg _410536_410536 ; 
   reg __410536_410536;
   reg _410537_410537 ; 
   reg __410537_410537;
   reg _410538_410538 ; 
   reg __410538_410538;
   reg _410539_410539 ; 
   reg __410539_410539;
   reg _410540_410540 ; 
   reg __410540_410540;
   reg _410541_410541 ; 
   reg __410541_410541;
   reg _410542_410542 ; 
   reg __410542_410542;
   reg _410543_410543 ; 
   reg __410543_410543;
   reg _410544_410544 ; 
   reg __410544_410544;
   reg _410545_410545 ; 
   reg __410545_410545;
   reg _410546_410546 ; 
   reg __410546_410546;
   reg _410547_410547 ; 
   reg __410547_410547;
   reg _410548_410548 ; 
   reg __410548_410548;
   reg _410549_410549 ; 
   reg __410549_410549;
   reg _410550_410550 ; 
   reg __410550_410550;
   reg _410551_410551 ; 
   reg __410551_410551;
   reg _410552_410552 ; 
   reg __410552_410552;
   reg _410553_410553 ; 
   reg __410553_410553;
   reg _410554_410554 ; 
   reg __410554_410554;
   reg _410555_410555 ; 
   reg __410555_410555;
   reg _410556_410556 ; 
   reg __410556_410556;
   reg _410557_410557 ; 
   reg __410557_410557;
   reg _410558_410558 ; 
   reg __410558_410558;
   reg _410559_410559 ; 
   reg __410559_410559;
   reg _410560_410560 ; 
   reg __410560_410560;
   reg _410561_410561 ; 
   reg __410561_410561;
   reg _410562_410562 ; 
   reg __410562_410562;
   reg _410563_410563 ; 
   reg __410563_410563;
   reg _410564_410564 ; 
   reg __410564_410564;
   reg _410565_410565 ; 
   reg __410565_410565;
   reg _410566_410566 ; 
   reg __410566_410566;
   reg _410567_410567 ; 
   reg __410567_410567;
   reg _410568_410568 ; 
   reg __410568_410568;
   reg _410569_410569 ; 
   reg __410569_410569;
   reg _410570_410570 ; 
   reg __410570_410570;
   reg _410571_410571 ; 
   reg __410571_410571;
   reg _410572_410572 ; 
   reg __410572_410572;
   reg _410573_410573 ; 
   reg __410573_410573;
   reg _410574_410574 ; 
   reg __410574_410574;
   reg _410575_410575 ; 
   reg __410575_410575;
   reg _410576_410576 ; 
   reg __410576_410576;
   reg _410577_410577 ; 
   reg __410577_410577;
   reg _410578_410578 ; 
   reg __410578_410578;
   reg _410579_410579 ; 
   reg __410579_410579;
   reg _410580_410580 ; 
   reg __410580_410580;
   reg _410581_410581 ; 
   reg __410581_410581;
   reg _410582_410582 ; 
   reg __410582_410582;
   reg _410583_410583 ; 
   reg __410583_410583;
   reg _410584_410584 ; 
   reg __410584_410584;
   reg _410585_410585 ; 
   reg __410585_410585;
   reg _410586_410586 ; 
   reg __410586_410586;
   reg _410587_410587 ; 
   reg __410587_410587;
   reg _410588_410588 ; 
   reg __410588_410588;
   reg _410589_410589 ; 
   reg __410589_410589;
   reg _410590_410590 ; 
   reg __410590_410590;
   reg _410591_410591 ; 
   reg __410591_410591;
   reg _410592_410592 ; 
   reg __410592_410592;
   reg _410593_410593 ; 
   reg __410593_410593;
   reg _410594_410594 ; 
   reg __410594_410594;
   reg _410595_410595 ; 
   reg __410595_410595;
   reg _410596_410596 ; 
   reg __410596_410596;
   reg _410597_410597 ; 
   reg __410597_410597;
   reg _410598_410598 ; 
   reg __410598_410598;
   reg _410599_410599 ; 
   reg __410599_410599;
   reg _410600_410600 ; 
   reg __410600_410600;
   reg _410601_410601 ; 
   reg __410601_410601;
   reg _410602_410602 ; 
   reg __410602_410602;
   reg _410603_410603 ; 
   reg __410603_410603;
   reg _410604_410604 ; 
   reg __410604_410604;
   reg _410605_410605 ; 
   reg __410605_410605;
   reg _410606_410606 ; 
   reg __410606_410606;
   reg _410607_410607 ; 
   reg __410607_410607;
   reg _410608_410608 ; 
   reg __410608_410608;
   reg _410609_410609 ; 
   reg __410609_410609;
   reg _410610_410610 ; 
   reg __410610_410610;
   reg _410611_410611 ; 
   reg __410611_410611;
   reg _410612_410612 ; 
   reg __410612_410612;
   reg _410613_410613 ; 
   reg __410613_410613;
   reg _410614_410614 ; 
   reg __410614_410614;
   reg _410615_410615 ; 
   reg __410615_410615;
   reg _410616_410616 ; 
   reg __410616_410616;
   reg _410617_410617 ; 
   reg __410617_410617;
   reg _410618_410618 ; 
   reg __410618_410618;
   reg _410619_410619 ; 
   reg __410619_410619;
   reg _410620_410620 ; 
   reg __410620_410620;
   reg _410621_410621 ; 
   reg __410621_410621;
   reg _410622_410622 ; 
   reg __410622_410622;
   reg _410623_410623 ; 
   reg __410623_410623;
   reg _410624_410624 ; 
   reg __410624_410624;
   reg _410625_410625 ; 
   reg __410625_410625;
   reg _410626_410626 ; 
   reg __410626_410626;
   reg _410627_410627 ; 
   reg __410627_410627;
   reg _410628_410628 ; 
   reg __410628_410628;
   reg _410629_410629 ; 
   reg __410629_410629;
   reg _410630_410630 ; 
   reg __410630_410630;
   reg _410631_410631 ; 
   reg __410631_410631;
   reg _410632_410632 ; 
   reg __410632_410632;
   reg _410633_410633 ; 
   reg __410633_410633;
   reg _410634_410634 ; 
   reg __410634_410634;
   reg _410635_410635 ; 
   reg __410635_410635;
   reg _410636_410636 ; 
   reg __410636_410636;
   reg _410637_410637 ; 
   reg __410637_410637;
   reg _410638_410638 ; 
   reg __410638_410638;
   reg _410639_410639 ; 
   reg __410639_410639;
   reg _410640_410640 ; 
   reg __410640_410640;
   reg _410641_410641 ; 
   reg __410641_410641;
   reg _410642_410642 ; 
   reg __410642_410642;
   reg _410643_410643 ; 
   reg __410643_410643;
   reg _410644_410644 ; 
   reg __410644_410644;
   reg _410645_410645 ; 
   reg __410645_410645;
   reg _410646_410646 ; 
   reg __410646_410646;
   reg _410647_410647 ; 
   reg __410647_410647;
   reg _410648_410648 ; 
   reg __410648_410648;
   reg _410649_410649 ; 
   reg __410649_410649;
   reg _410650_410650 ; 
   reg __410650_410650;
   reg _410651_410651 ; 
   reg __410651_410651;
   reg _410652_410652 ; 
   reg __410652_410652;
   reg _410653_410653 ; 
   reg __410653_410653;
   reg _410654_410654 ; 
   reg __410654_410654;
   reg _410655_410655 ; 
   reg __410655_410655;
   reg _410656_410656 ; 
   reg __410656_410656;
   reg _410657_410657 ; 
   reg __410657_410657;
   reg _410658_410658 ; 
   reg __410658_410658;
   reg _410659_410659 ; 
   reg __410659_410659;
   reg _410660_410660 ; 
   reg __410660_410660;
   reg _410661_410661 ; 
   reg __410661_410661;
   reg _410662_410662 ; 
   reg __410662_410662;
   reg _410663_410663 ; 
   reg __410663_410663;
   reg _410664_410664 ; 
   reg __410664_410664;
   reg _410665_410665 ; 
   reg __410665_410665;
   reg _410666_410666 ; 
   reg __410666_410666;
   reg _410667_410667 ; 
   reg __410667_410667;
   reg _410668_410668 ; 
   reg __410668_410668;
   reg _410669_410669 ; 
   reg __410669_410669;
   reg _410670_410670 ; 
   reg __410670_410670;
   reg _410671_410671 ; 
   reg __410671_410671;
   reg _410672_410672 ; 
   reg __410672_410672;
   reg _410673_410673 ; 
   reg __410673_410673;
   reg _410674_410674 ; 
   reg __410674_410674;
   reg _410675_410675 ; 
   reg __410675_410675;
   reg _410676_410676 ; 
   reg __410676_410676;
   reg _410677_410677 ; 
   reg __410677_410677;
   reg _410678_410678 ; 
   reg __410678_410678;
   reg _410679_410679 ; 
   reg __410679_410679;
   reg _410680_410680 ; 
   reg __410680_410680;
   reg _410681_410681 ; 
   reg __410681_410681;
   reg _410682_410682 ; 
   reg __410682_410682;
   reg _410683_410683 ; 
   reg __410683_410683;
   reg _410684_410684 ; 
   reg __410684_410684;
   reg _410685_410685 ; 
   reg __410685_410685;
   reg _410686_410686 ; 
   reg __410686_410686;
   reg _410687_410687 ; 
   reg __410687_410687;
   reg _410688_410688 ; 
   reg __410688_410688;
   reg _410689_410689 ; 
   reg __410689_410689;
   reg _410690_410690 ; 
   reg __410690_410690;
   reg _410691_410691 ; 
   reg __410691_410691;
   reg _410692_410692 ; 
   reg __410692_410692;
   reg _410693_410693 ; 
   reg __410693_410693;
   reg _410694_410694 ; 
   reg __410694_410694;
   reg _410695_410695 ; 
   reg __410695_410695;
   reg _410696_410696 ; 
   reg __410696_410696;
   reg _410697_410697 ; 
   reg __410697_410697;
   reg _410698_410698 ; 
   reg __410698_410698;
   reg _410699_410699 ; 
   reg __410699_410699;
   reg _410700_410700 ; 
   reg __410700_410700;
   reg _410701_410701 ; 
   reg __410701_410701;
   reg _410702_410702 ; 
   reg __410702_410702;
   reg _410703_410703 ; 
   reg __410703_410703;
   reg _410704_410704 ; 
   reg __410704_410704;
   reg _410705_410705 ; 
   reg __410705_410705;
   reg _410706_410706 ; 
   reg __410706_410706;
   reg _410707_410707 ; 
   reg __410707_410707;
   reg _410708_410708 ; 
   reg __410708_410708;
   reg _410709_410709 ; 
   reg __410709_410709;
   reg _410710_410710 ; 
   reg __410710_410710;
   reg _410711_410711 ; 
   reg __410711_410711;
   reg _410712_410712 ; 
   reg __410712_410712;
   reg _410713_410713 ; 
   reg __410713_410713;
   reg _410714_410714 ; 
   reg __410714_410714;
   reg _410715_410715 ; 
   reg __410715_410715;
   reg _410716_410716 ; 
   reg __410716_410716;
   reg _410717_410717 ; 
   reg __410717_410717;
   reg _410718_410718 ; 
   reg __410718_410718;
   reg _410719_410719 ; 
   reg __410719_410719;
   reg _410720_410720 ; 
   reg __410720_410720;
   reg _410721_410721 ; 
   reg __410721_410721;
   reg _410722_410722 ; 
   reg __410722_410722;
   reg _410723_410723 ; 
   reg __410723_410723;
   reg _410724_410724 ; 
   reg __410724_410724;
   reg _410725_410725 ; 
   reg __410725_410725;
   reg _410726_410726 ; 
   reg __410726_410726;
   reg _410727_410727 ; 
   reg __410727_410727;
   reg _410728_410728 ; 
   reg __410728_410728;
   reg _410729_410729 ; 
   reg __410729_410729;
   reg _410730_410730 ; 
   reg __410730_410730;
   reg _410731_410731 ; 
   reg __410731_410731;
   reg _410732_410732 ; 
   reg __410732_410732;
   reg _410733_410733 ; 
   reg __410733_410733;
   reg _410734_410734 ; 
   reg __410734_410734;
   reg _410735_410735 ; 
   reg __410735_410735;
   reg _410736_410736 ; 
   reg __410736_410736;
   reg _410737_410737 ; 
   reg __410737_410737;
   reg _410738_410738 ; 
   reg __410738_410738;
   reg _410739_410739 ; 
   reg __410739_410739;
   reg _410740_410740 ; 
   reg __410740_410740;
   reg _410741_410741 ; 
   reg __410741_410741;
   reg _410742_410742 ; 
   reg __410742_410742;
   reg _410743_410743 ; 
   reg __410743_410743;
   reg _410744_410744 ; 
   reg __410744_410744;
   reg _410745_410745 ; 
   reg __410745_410745;
   reg _410746_410746 ; 
   reg __410746_410746;
   reg _410747_410747 ; 
   reg __410747_410747;
   reg _410748_410748 ; 
   reg __410748_410748;
   reg _410749_410749 ; 
   reg __410749_410749;
   reg _410750_410750 ; 
   reg __410750_410750;
   reg _410751_410751 ; 
   reg __410751_410751;
   reg _410752_410752 ; 
   reg __410752_410752;
   reg _410753_410753 ; 
   reg __410753_410753;
   reg _410754_410754 ; 
   reg __410754_410754;
   reg _410755_410755 ; 
   reg __410755_410755;
   reg _410756_410756 ; 
   reg __410756_410756;
   reg _410757_410757 ; 
   reg __410757_410757;
   reg _410758_410758 ; 
   reg __410758_410758;
   reg _410759_410759 ; 
   reg __410759_410759;
   reg _410760_410760 ; 
   reg __410760_410760;
   reg _410761_410761 ; 
   reg __410761_410761;
   reg _410762_410762 ; 
   reg __410762_410762;
   reg _410763_410763 ; 
   reg __410763_410763;
   reg _410764_410764 ; 
   reg __410764_410764;
   reg _410765_410765 ; 
   reg __410765_410765;
   reg _410766_410766 ; 
   reg __410766_410766;
   reg _410767_410767 ; 
   reg __410767_410767;
   reg _410768_410768 ; 
   reg __410768_410768;
   reg _410769_410769 ; 
   reg __410769_410769;
   reg _410770_410770 ; 
   reg __410770_410770;
   reg _410771_410771 ; 
   reg __410771_410771;
   reg _410772_410772 ; 
   reg __410772_410772;
   reg _410773_410773 ; 
   reg __410773_410773;
   reg _410774_410774 ; 
   reg __410774_410774;
   reg _410775_410775 ; 
   reg __410775_410775;
   reg _410776_410776 ; 
   reg __410776_410776;
   reg _410777_410777 ; 
   reg __410777_410777;
   reg _410778_410778 ; 
   reg __410778_410778;
   reg _410779_410779 ; 
   reg __410779_410779;
   reg _410780_410780 ; 
   reg __410780_410780;
   reg _410781_410781 ; 
   reg __410781_410781;
   reg _410782_410782 ; 
   reg __410782_410782;
   reg _410783_410783 ; 
   reg __410783_410783;
   reg _410784_410784 ; 
   reg __410784_410784;
   reg _410785_410785 ; 
   reg __410785_410785;
   reg _410786_410786 ; 
   reg __410786_410786;
   reg _410787_410787 ; 
   reg __410787_410787;
   reg _410788_410788 ; 
   reg __410788_410788;
   reg _410789_410789 ; 
   reg __410789_410789;
   reg _410790_410790 ; 
   reg __410790_410790;
   reg _410791_410791 ; 
   reg __410791_410791;
   reg _410792_410792 ; 
   reg __410792_410792;
   reg _410793_410793 ; 
   reg __410793_410793;
   reg _410794_410794 ; 
   reg __410794_410794;
   reg _410795_410795 ; 
   reg __410795_410795;
   reg _410796_410796 ; 
   reg __410796_410796;
   reg _410797_410797 ; 
   reg __410797_410797;
   reg _410798_410798 ; 
   reg __410798_410798;
   reg _410799_410799 ; 
   reg __410799_410799;
   reg _410800_410800 ; 
   reg __410800_410800;
   reg _410801_410801 ; 
   reg __410801_410801;
   reg _410802_410802 ; 
   reg __410802_410802;
   reg _410803_410803 ; 
   reg __410803_410803;
   reg _410804_410804 ; 
   reg __410804_410804;
   reg _410805_410805 ; 
   reg __410805_410805;
   reg _410806_410806 ; 
   reg __410806_410806;
   reg _410807_410807 ; 
   reg __410807_410807;
   reg _410808_410808 ; 
   reg __410808_410808;
   reg _410809_410809 ; 
   reg __410809_410809;
   reg _410810_410810 ; 
   reg __410810_410810;
   reg _410811_410811 ; 
   reg __410811_410811;
   reg _410812_410812 ; 
   reg __410812_410812;
   reg _410813_410813 ; 
   reg __410813_410813;
   reg _410814_410814 ; 
   reg __410814_410814;
   reg _410815_410815 ; 
   reg __410815_410815;
   reg _410816_410816 ; 
   reg __410816_410816;
   reg _410817_410817 ; 
   reg __410817_410817;
   reg _410818_410818 ; 
   reg __410818_410818;
   reg _410819_410819 ; 
   reg __410819_410819;
   reg _410820_410820 ; 
   reg __410820_410820;
   reg _410821_410821 ; 
   reg __410821_410821;
   reg _410822_410822 ; 
   reg __410822_410822;
   reg _410823_410823 ; 
   reg __410823_410823;
   reg _410824_410824 ; 
   reg __410824_410824;
   reg _410825_410825 ; 
   reg __410825_410825;
   reg _410826_410826 ; 
   reg __410826_410826;
   reg _410827_410827 ; 
   reg __410827_410827;
   reg _410828_410828 ; 
   reg __410828_410828;
   reg _410829_410829 ; 
   reg __410829_410829;
   reg _410830_410830 ; 
   reg __410830_410830;
   reg _410831_410831 ; 
   reg __410831_410831;
   reg _410832_410832 ; 
   reg __410832_410832;
   reg _410833_410833 ; 
   reg __410833_410833;
   reg _410834_410834 ; 
   reg __410834_410834;
   reg _410835_410835 ; 
   reg __410835_410835;
   reg _410836_410836 ; 
   reg __410836_410836;
   reg _410837_410837 ; 
   reg __410837_410837;
   reg _410838_410838 ; 
   reg __410838_410838;
   reg _410839_410839 ; 
   reg __410839_410839;
   reg _410840_410840 ; 
   reg __410840_410840;
   reg _410841_410841 ; 
   reg __410841_410841;
   reg _410842_410842 ; 
   reg __410842_410842;
   reg _410843_410843 ; 
   reg __410843_410843;
   reg _410844_410844 ; 
   reg __410844_410844;
   reg _410845_410845 ; 
   reg __410845_410845;
   reg _410846_410846 ; 
   reg __410846_410846;
   reg _410847_410847 ; 
   reg __410847_410847;
   reg _410848_410848 ; 
   reg __410848_410848;
   reg _410849_410849 ; 
   reg __410849_410849;
   reg _410850_410850 ; 
   reg __410850_410850;
   reg _410851_410851 ; 
   reg __410851_410851;
   reg _410852_410852 ; 
   reg __410852_410852;
   reg _410853_410853 ; 
   reg __410853_410853;
   reg _410854_410854 ; 
   reg __410854_410854;
   reg _410855_410855 ; 
   reg __410855_410855;
   reg _410856_410856 ; 
   reg __410856_410856;
   reg _410857_410857 ; 
   reg __410857_410857;
   reg _410858_410858 ; 
   reg __410858_410858;
   reg _410859_410859 ; 
   reg __410859_410859;
   reg _410860_410860 ; 
   reg __410860_410860;
   reg _410861_410861 ; 
   reg __410861_410861;
   reg _410862_410862 ; 
   reg __410862_410862;
   reg _410863_410863 ; 
   reg __410863_410863;
   reg _410864_410864 ; 
   reg __410864_410864;
   reg _410865_410865 ; 
   reg __410865_410865;
   reg _410866_410866 ; 
   reg __410866_410866;
   reg _410867_410867 ; 
   reg __410867_410867;
   reg _410868_410868 ; 
   reg __410868_410868;
   reg _410869_410869 ; 
   reg __410869_410869;
   reg _410870_410870 ; 
   reg __410870_410870;
   reg _410871_410871 ; 
   reg __410871_410871;
   reg _410872_410872 ; 
   reg __410872_410872;
   reg _410873_410873 ; 
   reg __410873_410873;
   reg _410874_410874 ; 
   reg __410874_410874;
   reg _410875_410875 ; 
   reg __410875_410875;
   reg _410876_410876 ; 
   reg __410876_410876;
   reg _410877_410877 ; 
   reg __410877_410877;
   reg _410878_410878 ; 
   reg __410878_410878;
   reg _410879_410879 ; 
   reg __410879_410879;
   reg _410880_410880 ; 
   reg __410880_410880;
   reg _410881_410881 ; 
   reg __410881_410881;
   reg _410882_410882 ; 
   reg __410882_410882;
   reg _410883_410883 ; 
   reg __410883_410883;
   reg _410884_410884 ; 
   reg __410884_410884;
   reg _410885_410885 ; 
   reg __410885_410885;
   reg _410886_410886 ; 
   reg __410886_410886;
   reg _410887_410887 ; 
   reg __410887_410887;
   reg _410888_410888 ; 
   reg __410888_410888;
   reg _410889_410889 ; 
   reg __410889_410889;
   reg _410890_410890 ; 
   reg __410890_410890;
   reg _410891_410891 ; 
   reg __410891_410891;
   reg _410892_410892 ; 
   reg __410892_410892;
   reg _410893_410893 ; 
   reg __410893_410893;
   reg _410894_410894 ; 
   reg __410894_410894;
   reg _410895_410895 ; 
   reg __410895_410895;
   reg _410896_410896 ; 
   reg __410896_410896;
   reg _410897_410897 ; 
   reg __410897_410897;
   reg _410898_410898 ; 
   reg __410898_410898;
   reg _410899_410899 ; 
   reg __410899_410899;
   reg _410900_410900 ; 
   reg __410900_410900;
   reg _410901_410901 ; 
   reg __410901_410901;
   reg _410902_410902 ; 
   reg __410902_410902;
   reg _410903_410903 ; 
   reg __410903_410903;
   reg _410904_410904 ; 
   reg __410904_410904;
   reg _410905_410905 ; 
   reg __410905_410905;
   reg _410906_410906 ; 
   reg __410906_410906;
   reg _410907_410907 ; 
   reg __410907_410907;
   reg _410908_410908 ; 
   reg __410908_410908;
   reg _410909_410909 ; 
   reg __410909_410909;
   reg _410910_410910 ; 
   reg __410910_410910;
   reg _410911_410911 ; 
   reg __410911_410911;
   reg _410912_410912 ; 
   reg __410912_410912;
   reg _410913_410913 ; 
   reg __410913_410913;
   reg _410914_410914 ; 
   reg __410914_410914;
   reg _410915_410915 ; 
   reg __410915_410915;
   reg _410916_410916 ; 
   reg __410916_410916;
   reg _410917_410917 ; 
   reg __410917_410917;
   reg _410918_410918 ; 
   reg __410918_410918;
   reg _410919_410919 ; 
   reg __410919_410919;
   reg _410920_410920 ; 
   reg __410920_410920;
   reg _410921_410921 ; 
   reg __410921_410921;
   reg _410922_410922 ; 
   reg __410922_410922;
   reg _410923_410923 ; 
   reg __410923_410923;
   reg _410924_410924 ; 
   reg __410924_410924;
   reg _410925_410925 ; 
   reg __410925_410925;
   reg _410926_410926 ; 
   reg __410926_410926;
   reg _410927_410927 ; 
   reg __410927_410927;
   reg _410928_410928 ; 
   reg __410928_410928;
   reg _410929_410929 ; 
   reg __410929_410929;
   reg _410930_410930 ; 
   reg __410930_410930;
   reg _410931_410931 ; 
   reg __410931_410931;
   reg _410932_410932 ; 
   reg __410932_410932;
   reg _410933_410933 ; 
   reg __410933_410933;
   reg _410934_410934 ; 
   reg __410934_410934;
   reg _410935_410935 ; 
   reg __410935_410935;
   reg _410936_410936 ; 
   reg __410936_410936;
   reg _410937_410937 ; 
   reg __410937_410937;
   reg _410938_410938 ; 
   reg __410938_410938;
   reg _410939_410939 ; 
   reg __410939_410939;
   reg _410940_410940 ; 
   reg __410940_410940;
   reg _410941_410941 ; 
   reg __410941_410941;
   reg _410942_410942 ; 
   reg __410942_410942;
   reg _410943_410943 ; 
   reg __410943_410943;
   reg _410944_410944 ; 
   reg __410944_410944;
   reg _410945_410945 ; 
   reg __410945_410945;
   reg _410946_410946 ; 
   reg __410946_410946;
   reg _410947_410947 ; 
   reg __410947_410947;
   reg _410948_410948 ; 
   reg __410948_410948;
   reg _410949_410949 ; 
   reg __410949_410949;
   reg _410950_410950 ; 
   reg __410950_410950;
   reg _410951_410951 ; 
   reg __410951_410951;
   reg _410952_410952 ; 
   reg __410952_410952;
   reg _410953_410953 ; 
   reg __410953_410953;
   reg _410954_410954 ; 
   reg __410954_410954;
   reg _410955_410955 ; 
   reg __410955_410955;
   reg _410956_410956 ; 
   reg __410956_410956;
   reg _410957_410957 ; 
   reg __410957_410957;
   reg _410958_410958 ; 
   reg __410958_410958;
   reg _410959_410959 ; 
   reg __410959_410959;
   reg _410960_410960 ; 
   reg __410960_410960;
   reg _410961_410961 ; 
   reg __410961_410961;
   reg _410962_410962 ; 
   reg __410962_410962;
   reg _410963_410963 ; 
   reg __410963_410963;
   reg _410964_410964 ; 
   reg __410964_410964;
   reg _410965_410965 ; 
   reg __410965_410965;
   reg _410966_410966 ; 
   reg __410966_410966;
   reg _410967_410967 ; 
   reg __410967_410967;
   reg _410968_410968 ; 
   reg __410968_410968;
   reg _410969_410969 ; 
   reg __410969_410969;
   reg _410970_410970 ; 
   reg __410970_410970;
   reg _410971_410971 ; 
   reg __410971_410971;
   reg _410972_410972 ; 
   reg __410972_410972;
   reg _410973_410973 ; 
   reg __410973_410973;
   reg _410974_410974 ; 
   reg __410974_410974;
   reg _410975_410975 ; 
   reg __410975_410975;
   reg _410976_410976 ; 
   reg __410976_410976;
   reg _410977_410977 ; 
   reg __410977_410977;
   reg _410978_410978 ; 
   reg __410978_410978;
   reg _410979_410979 ; 
   reg __410979_410979;
   reg _410980_410980 ; 
   reg __410980_410980;
   reg _410981_410981 ; 
   reg __410981_410981;
   reg _410982_410982 ; 
   reg __410982_410982;
   reg _410983_410983 ; 
   reg __410983_410983;
   reg _410984_410984 ; 
   reg __410984_410984;
   reg _410985_410985 ; 
   reg __410985_410985;
   reg _410986_410986 ; 
   reg __410986_410986;
   reg _410987_410987 ; 
   reg __410987_410987;
   reg _410988_410988 ; 
   reg __410988_410988;
   reg _410989_410989 ; 
   reg __410989_410989;
   reg _410990_410990 ; 
   reg __410990_410990;
   reg _410991_410991 ; 
   reg __410991_410991;
   reg _410992_410992 ; 
   reg __410992_410992;
   reg _410993_410993 ; 
   reg __410993_410993;
   reg _410994_410994 ; 
   reg __410994_410994;
   reg _410995_410995 ; 
   reg __410995_410995;
   reg _410996_410996 ; 
   reg __410996_410996;
   reg _410997_410997 ; 
   reg __410997_410997;
   reg _410998_410998 ; 
   reg __410998_410998;
   reg _410999_410999 ; 
   reg __410999_410999;
   reg _411000_411000 ; 
   reg __411000_411000;
   reg _411001_411001 ; 
   reg __411001_411001;
   reg _411002_411002 ; 
   reg __411002_411002;
   reg _411003_411003 ; 
   reg __411003_411003;
   reg _411004_411004 ; 
   reg __411004_411004;
   reg _411005_411005 ; 
   reg __411005_411005;
   reg _411006_411006 ; 
   reg __411006_411006;
   reg _411007_411007 ; 
   reg __411007_411007;
   reg _411008_411008 ; 
   reg __411008_411008;
   reg _411009_411009 ; 
   reg __411009_411009;
   reg _411010_411010 ; 
   reg __411010_411010;
   reg _411011_411011 ; 
   reg __411011_411011;
   reg _411012_411012 ; 
   reg __411012_411012;
   reg _411013_411013 ; 
   reg __411013_411013;
   reg _411014_411014 ; 
   reg __411014_411014;
   reg _411015_411015 ; 
   reg __411015_411015;
   reg _411016_411016 ; 
   reg __411016_411016;
   reg _411017_411017 ; 
   reg __411017_411017;
   reg _411018_411018 ; 
   reg __411018_411018;
   reg _411019_411019 ; 
   reg __411019_411019;
   reg _411020_411020 ; 
   reg __411020_411020;
   reg _411021_411021 ; 
   reg __411021_411021;
   reg _411022_411022 ; 
   reg __411022_411022;
   reg _411023_411023 ; 
   reg __411023_411023;
   reg _411024_411024 ; 
   reg __411024_411024;
   reg _411025_411025 ; 
   reg __411025_411025;
   reg _411026_411026 ; 
   reg __411026_411026;
   reg _411027_411027 ; 
   reg __411027_411027;
   reg _411028_411028 ; 
   reg __411028_411028;
   reg _411029_411029 ; 
   reg __411029_411029;
   reg _411030_411030 ; 
   reg __411030_411030;
   reg _411031_411031 ; 
   reg __411031_411031;
   reg _411032_411032 ; 
   reg __411032_411032;
   reg _411033_411033 ; 
   reg __411033_411033;
   reg _411034_411034 ; 
   reg __411034_411034;
   reg _411035_411035 ; 
   reg __411035_411035;
   reg _411036_411036 ; 
   reg __411036_411036;
   reg _411037_411037 ; 
   reg __411037_411037;
   reg _411038_411038 ; 
   reg __411038_411038;
   reg _411039_411039 ; 
   reg __411039_411039;
   reg _411040_411040 ; 
   reg __411040_411040;
   reg _411041_411041 ; 
   reg __411041_411041;
   reg _411042_411042 ; 
   reg __411042_411042;
   reg _411043_411043 ; 
   reg __411043_411043;
   reg _411044_411044 ; 
   reg __411044_411044;
   reg _411045_411045 ; 
   reg __411045_411045;
   reg _411046_411046 ; 
   reg __411046_411046;
   reg _411047_411047 ; 
   reg __411047_411047;
   reg _411048_411048 ; 
   reg __411048_411048;
   reg _411049_411049 ; 
   reg __411049_411049;
   reg _411050_411050 ; 
   reg __411050_411050;
   reg _411051_411051 ; 
   reg __411051_411051;
   reg _411052_411052 ; 
   reg __411052_411052;
   reg _411053_411053 ; 
   reg __411053_411053;
   reg _411054_411054 ; 
   reg __411054_411054;
   reg _411055_411055 ; 
   reg __411055_411055;
   reg _411056_411056 ; 
   reg __411056_411056;
   reg _411057_411057 ; 
   reg __411057_411057;
   reg _411058_411058 ; 
   reg __411058_411058;
   reg _411059_411059 ; 
   reg __411059_411059;
   reg _411060_411060 ; 
   reg __411060_411060;
   reg _411061_411061 ; 
   reg __411061_411061;
   reg _411062_411062 ; 
   reg __411062_411062;
   reg _411063_411063 ; 
   reg __411063_411063;
   reg _411064_411064 ; 
   reg __411064_411064;
   reg _411065_411065 ; 
   reg __411065_411065;
   reg _411066_411066 ; 
   reg __411066_411066;
   reg _411067_411067 ; 
   reg __411067_411067;
   reg _411068_411068 ; 
   reg __411068_411068;
   reg _411069_411069 ; 
   reg __411069_411069;
   reg _411070_411070 ; 
   reg __411070_411070;
   reg _411071_411071 ; 
   reg __411071_411071;
   reg _411072_411072 ; 
   reg __411072_411072;
   reg _411073_411073 ; 
   reg __411073_411073;
   reg _411074_411074 ; 
   reg __411074_411074;
   reg _411075_411075 ; 
   reg __411075_411075;
   reg _411076_411076 ; 
   reg __411076_411076;
   reg _411077_411077 ; 
   reg __411077_411077;
   reg _411078_411078 ; 
   reg __411078_411078;
   reg _411079_411079 ; 
   reg __411079_411079;
   reg _411080_411080 ; 
   reg __411080_411080;
   reg _411081_411081 ; 
   reg __411081_411081;
   reg _411082_411082 ; 
   reg __411082_411082;
   reg _411083_411083 ; 
   reg __411083_411083;
   reg _411084_411084 ; 
   reg __411084_411084;
   reg _411085_411085 ; 
   reg __411085_411085;
   reg _411086_411086 ; 
   reg __411086_411086;
   reg _411087_411087 ; 
   reg __411087_411087;
   reg _411088_411088 ; 
   reg __411088_411088;
   reg _411089_411089 ; 
   reg __411089_411089;
   reg _411090_411090 ; 
   reg __411090_411090;
   reg _411091_411091 ; 
   reg __411091_411091;
   reg _411092_411092 ; 
   reg __411092_411092;
   reg _411093_411093 ; 
   reg __411093_411093;
   reg _411094_411094 ; 
   reg __411094_411094;
   reg _411095_411095 ; 
   reg __411095_411095;
   reg _411096_411096 ; 
   reg __411096_411096;
   reg _411097_411097 ; 
   reg __411097_411097;
   reg _411098_411098 ; 
   reg __411098_411098;
   reg _411099_411099 ; 
   reg __411099_411099;
   reg _411100_411100 ; 
   reg __411100_411100;
   reg _411101_411101 ; 
   reg __411101_411101;
   reg _411102_411102 ; 
   reg __411102_411102;
   reg _411103_411103 ; 
   reg __411103_411103;
   reg _411104_411104 ; 
   reg __411104_411104;
   reg _411105_411105 ; 
   reg __411105_411105;
   reg _411106_411106 ; 
   reg __411106_411106;
   reg _411107_411107 ; 
   reg __411107_411107;
   reg _411108_411108 ; 
   reg __411108_411108;
   reg _411109_411109 ; 
   reg __411109_411109;
   reg _411110_411110 ; 
   reg __411110_411110;
   reg _411111_411111 ; 
   reg __411111_411111;
   reg _411112_411112 ; 
   reg __411112_411112;
   reg _411113_411113 ; 
   reg __411113_411113;
   reg _411114_411114 ; 
   reg __411114_411114;
   reg _411115_411115 ; 
   reg __411115_411115;
   reg _411116_411116 ; 
   reg __411116_411116;
   reg _411117_411117 ; 
   reg __411117_411117;
   reg _411118_411118 ; 
   reg __411118_411118;
   reg _411119_411119 ; 
   reg __411119_411119;
   reg _411120_411120 ; 
   reg __411120_411120;
   reg _411121_411121 ; 
   reg __411121_411121;
   reg _411122_411122 ; 
   reg __411122_411122;
   reg _411123_411123 ; 
   reg __411123_411123;
   reg _411124_411124 ; 
   reg __411124_411124;
   reg _411125_411125 ; 
   reg __411125_411125;
   reg _411126_411126 ; 
   reg __411126_411126;
   reg _411127_411127 ; 
   reg __411127_411127;
   reg _411128_411128 ; 
   reg __411128_411128;
   reg _411129_411129 ; 
   reg __411129_411129;
   reg _411130_411130 ; 
   reg __411130_411130;
   reg _411131_411131 ; 
   reg __411131_411131;
   reg _411132_411132 ; 
   reg __411132_411132;
   reg _411133_411133 ; 
   reg __411133_411133;
   reg _411134_411134 ; 
   reg __411134_411134;
   reg _411135_411135 ; 
   reg __411135_411135;
   reg _411136_411136 ; 
   reg __411136_411136;
   reg _411137_411137 ; 
   reg __411137_411137;
   reg _411138_411138 ; 
   reg __411138_411138;
   reg _411139_411139 ; 
   reg __411139_411139;
   reg _411140_411140 ; 
   reg __411140_411140;
   reg _411141_411141 ; 
   reg __411141_411141;
   reg _411142_411142 ; 
   reg __411142_411142;
   reg _411143_411143 ; 
   reg __411143_411143;
   reg _411144_411144 ; 
   reg __411144_411144;
   reg _411145_411145 ; 
   reg __411145_411145;
   reg _411146_411146 ; 
   reg __411146_411146;
   reg _411147_411147 ; 
   reg __411147_411147;
   reg _411148_411148 ; 
   reg __411148_411148;
   reg _411149_411149 ; 
   reg __411149_411149;
   reg _411150_411150 ; 
   reg __411150_411150;
   reg _411151_411151 ; 
   reg __411151_411151;
   reg _411152_411152 ; 
   reg __411152_411152;
   reg _411153_411153 ; 
   reg __411153_411153;
   reg _411154_411154 ; 
   reg __411154_411154;
   reg _411155_411155 ; 
   reg __411155_411155;
   reg _411156_411156 ; 
   reg __411156_411156;
   reg _411157_411157 ; 
   reg __411157_411157;
   reg _411158_411158 ; 
   reg __411158_411158;
   reg _411159_411159 ; 
   reg __411159_411159;
   reg _411160_411160 ; 
   reg __411160_411160;
   reg _411161_411161 ; 
   reg __411161_411161;
   reg _411162_411162 ; 
   reg __411162_411162;
   reg _411163_411163 ; 
   reg __411163_411163;
   reg _411164_411164 ; 
   reg __411164_411164;
   reg _411165_411165 ; 
   reg __411165_411165;
   reg _411166_411166 ; 
   reg __411166_411166;
   reg _411167_411167 ; 
   reg __411167_411167;
   reg _411168_411168 ; 
   reg __411168_411168;
   reg _411169_411169 ; 
   reg __411169_411169;
   reg _411170_411170 ; 
   reg __411170_411170;
   reg _411171_411171 ; 
   reg __411171_411171;
   reg _411172_411172 ; 
   reg __411172_411172;
   reg _411173_411173 ; 
   reg __411173_411173;
   reg _411174_411174 ; 
   reg __411174_411174;
   reg _411175_411175 ; 
   reg __411175_411175;
   reg _411176_411176 ; 
   reg __411176_411176;
   reg _411177_411177 ; 
   reg __411177_411177;
   reg _411178_411178 ; 
   reg __411178_411178;
   reg _411179_411179 ; 
   reg __411179_411179;
   reg _411180_411180 ; 
   reg __411180_411180;
   reg _411181_411181 ; 
   reg __411181_411181;
   reg _411182_411182 ; 
   reg __411182_411182;
   reg _411183_411183 ; 
   reg __411183_411183;
   reg _411184_411184 ; 
   reg __411184_411184;
   reg _411185_411185 ; 
   reg __411185_411185;
   reg _411186_411186 ; 
   reg __411186_411186;
   reg _411187_411187 ; 
   reg __411187_411187;
   reg _411188_411188 ; 
   reg __411188_411188;
   reg _411189_411189 ; 
   reg __411189_411189;
   reg _411190_411190 ; 
   reg __411190_411190;
   reg _411191_411191 ; 
   reg __411191_411191;
   reg _411192_411192 ; 
   reg __411192_411192;
   reg _411193_411193 ; 
   reg __411193_411193;
   reg _411194_411194 ; 
   reg __411194_411194;
   reg _411195_411195 ; 
   reg __411195_411195;
   reg _411196_411196 ; 
   reg __411196_411196;
   reg _411197_411197 ; 
   reg __411197_411197;
   reg _411198_411198 ; 
   reg __411198_411198;
   reg _411199_411199 ; 
   reg __411199_411199;
   reg _411200_411200 ; 
   reg __411200_411200;
   reg _411201_411201 ; 
   reg __411201_411201;
   reg _411202_411202 ; 
   reg __411202_411202;
   reg _411203_411203 ; 
   reg __411203_411203;
   reg _411204_411204 ; 
   reg __411204_411204;
   reg _411205_411205 ; 
   reg __411205_411205;
   reg _411206_411206 ; 
   reg __411206_411206;
   reg _411207_411207 ; 
   reg __411207_411207;
   reg _411208_411208 ; 
   reg __411208_411208;
   reg _411209_411209 ; 
   reg __411209_411209;
   reg _411210_411210 ; 
   reg __411210_411210;
   reg _411211_411211 ; 
   reg __411211_411211;
   reg _411212_411212 ; 
   reg __411212_411212;
   reg _411213_411213 ; 
   reg __411213_411213;
   reg _411214_411214 ; 
   reg __411214_411214;
   reg _411215_411215 ; 
   reg __411215_411215;
   reg _411216_411216 ; 
   reg __411216_411216;
   reg _411217_411217 ; 
   reg __411217_411217;
   reg _411218_411218 ; 
   reg __411218_411218;
   reg _411219_411219 ; 
   reg __411219_411219;
   reg _411220_411220 ; 
   reg __411220_411220;
   reg _411221_411221 ; 
   reg __411221_411221;
   reg _411222_411222 ; 
   reg __411222_411222;
   reg _411223_411223 ; 
   reg __411223_411223;
   reg _411224_411224 ; 
   reg __411224_411224;
   reg _411225_411225 ; 
   reg __411225_411225;
   reg _411226_411226 ; 
   reg __411226_411226;
   reg _411227_411227 ; 
   reg __411227_411227;
   reg _411228_411228 ; 
   reg __411228_411228;
   reg _411229_411229 ; 
   reg __411229_411229;
   reg _411230_411230 ; 
   reg __411230_411230;
   reg _411231_411231 ; 
   reg __411231_411231;
   reg _411232_411232 ; 
   reg __411232_411232;
   reg _411233_411233 ; 
   reg __411233_411233;
   reg _411234_411234 ; 
   reg __411234_411234;
   reg _411235_411235 ; 
   reg __411235_411235;
   reg _411236_411236 ; 
   reg __411236_411236;
   reg _411237_411237 ; 
   reg __411237_411237;
   reg _411238_411238 ; 
   reg __411238_411238;
   reg _411239_411239 ; 
   reg __411239_411239;
   reg _411240_411240 ; 
   reg __411240_411240;
   reg _411241_411241 ; 
   reg __411241_411241;
   reg _411242_411242 ; 
   reg __411242_411242;
   reg _411243_411243 ; 
   reg __411243_411243;
   reg _411244_411244 ; 
   reg __411244_411244;
   reg _411245_411245 ; 
   reg __411245_411245;
   reg _411246_411246 ; 
   reg __411246_411246;
   reg _411247_411247 ; 
   reg __411247_411247;
   reg _411248_411248 ; 
   reg __411248_411248;
   reg _411249_411249 ; 
   reg __411249_411249;
   reg _411250_411250 ; 
   reg __411250_411250;
   reg _411251_411251 ; 
   reg __411251_411251;
   reg _411252_411252 ; 
   reg __411252_411252;
   reg _411253_411253 ; 
   reg __411253_411253;
   reg _411254_411254 ; 
   reg __411254_411254;
   reg _411255_411255 ; 
   reg __411255_411255;
   reg _411256_411256 ; 
   reg __411256_411256;
   reg _411257_411257 ; 
   reg __411257_411257;
   reg _411258_411258 ; 
   reg __411258_411258;
   reg _411259_411259 ; 
   reg __411259_411259;
   reg _411260_411260 ; 
   reg __411260_411260;
   reg _411261_411261 ; 
   reg __411261_411261;
   reg _411262_411262 ; 
   reg __411262_411262;
   reg _411263_411263 ; 
   reg __411263_411263;
   reg _411264_411264 ; 
   reg __411264_411264;
   reg _411265_411265 ; 
   reg __411265_411265;
   reg _411266_411266 ; 
   reg __411266_411266;
   reg _411267_411267 ; 
   reg __411267_411267;
   reg _411268_411268 ; 
   reg __411268_411268;
   reg _411269_411269 ; 
   reg __411269_411269;
   reg _411270_411270 ; 
   reg __411270_411270;
   reg _411271_411271 ; 
   reg __411271_411271;
   reg _411272_411272 ; 
   reg __411272_411272;
   reg _411273_411273 ; 
   reg __411273_411273;
   reg _411274_411274 ; 
   reg __411274_411274;
   reg _411275_411275 ; 
   reg __411275_411275;
   reg _411276_411276 ; 
   reg __411276_411276;
   reg _411277_411277 ; 
   reg __411277_411277;
   reg _411278_411278 ; 
   reg __411278_411278;
   reg _411279_411279 ; 
   reg __411279_411279;
   reg _411280_411280 ; 
   reg __411280_411280;
   reg _411281_411281 ; 
   reg __411281_411281;
   reg _411282_411282 ; 
   reg __411282_411282;
   reg _411283_411283 ; 
   reg __411283_411283;
   reg _411284_411284 ; 
   reg __411284_411284;
   reg _411285_411285 ; 
   reg __411285_411285;
   reg _411286_411286 ; 
   reg __411286_411286;
   reg _411287_411287 ; 
   reg __411287_411287;
   reg _411288_411288 ; 
   reg __411288_411288;
   reg _411289_411289 ; 
   reg __411289_411289;
   reg _411290_411290 ; 
   reg __411290_411290;
   reg _411291_411291 ; 
   reg __411291_411291;
   reg _411292_411292 ; 
   reg __411292_411292;
   reg _411293_411293 ; 
   reg __411293_411293;
   reg _411294_411294 ; 
   reg __411294_411294;
   reg _411295_411295 ; 
   reg __411295_411295;
   reg _411296_411296 ; 
   reg __411296_411296;
   reg _411297_411297 ; 
   reg __411297_411297;
   reg _411298_411298 ; 
   reg __411298_411298;
   reg _411299_411299 ; 
   reg __411299_411299;
   reg _411300_411300 ; 
   reg __411300_411300;
   reg _411301_411301 ; 
   reg __411301_411301;
   reg _411302_411302 ; 
   reg __411302_411302;
   reg _411303_411303 ; 
   reg __411303_411303;
   reg _411304_411304 ; 
   reg __411304_411304;
   reg _411305_411305 ; 
   reg __411305_411305;
   reg _411306_411306 ; 
   reg __411306_411306;
   reg _411307_411307 ; 
   reg __411307_411307;
   reg _411308_411308 ; 
   reg __411308_411308;
   reg _411309_411309 ; 
   reg __411309_411309;
   reg _411310_411310 ; 
   reg __411310_411310;
   reg _411311_411311 ; 
   reg __411311_411311;
   reg _411312_411312 ; 
   reg __411312_411312;
   reg _411313_411313 ; 
   reg __411313_411313;
   reg _411314_411314 ; 
   reg __411314_411314;
   reg _411315_411315 ; 
   reg __411315_411315;
   reg _411316_411316 ; 
   reg __411316_411316;
   reg _411317_411317 ; 
   reg __411317_411317;
   reg _411318_411318 ; 
   reg __411318_411318;
   reg _411319_411319 ; 
   reg __411319_411319;
   reg _411320_411320 ; 
   reg __411320_411320;
   reg _411321_411321 ; 
   reg __411321_411321;
   reg _411322_411322 ; 
   reg __411322_411322;
   reg _411323_411323 ; 
   reg __411323_411323;
   reg _411324_411324 ; 
   reg __411324_411324;
   reg _411325_411325 ; 
   reg __411325_411325;
   reg _411326_411326 ; 
   reg __411326_411326;
   reg _411327_411327 ; 
   reg __411327_411327;
   reg _411328_411328 ; 
   reg __411328_411328;
   reg _411329_411329 ; 
   reg __411329_411329;
   reg _411330_411330 ; 
   reg __411330_411330;
   reg _411331_411331 ; 
   reg __411331_411331;
   reg _411332_411332 ; 
   reg __411332_411332;
   reg _411333_411333 ; 
   reg __411333_411333;
   reg _411334_411334 ; 
   reg __411334_411334;
   reg _411335_411335 ; 
   reg __411335_411335;
   reg _411336_411336 ; 
   reg __411336_411336;
   reg _411337_411337 ; 
   reg __411337_411337;
   reg _411338_411338 ; 
   reg __411338_411338;
   reg _411339_411339 ; 
   reg __411339_411339;
   reg _411340_411340 ; 
   reg __411340_411340;
   reg _411341_411341 ; 
   reg __411341_411341;
   reg _411342_411342 ; 
   reg __411342_411342;
   reg _411343_411343 ; 
   reg __411343_411343;
   reg _411344_411344 ; 
   reg __411344_411344;
   reg _411345_411345 ; 
   reg __411345_411345;
   reg _411346_411346 ; 
   reg __411346_411346;
   reg _411347_411347 ; 
   reg __411347_411347;
   reg _411348_411348 ; 
   reg __411348_411348;
   reg _411349_411349 ; 
   reg __411349_411349;
   reg _411350_411350 ; 
   reg __411350_411350;
   reg _411351_411351 ; 
   reg __411351_411351;
   reg _411352_411352 ; 
   reg __411352_411352;
   reg _411353_411353 ; 
   reg __411353_411353;
   reg _411354_411354 ; 
   reg __411354_411354;
   reg _411355_411355 ; 
   reg __411355_411355;
   reg _411356_411356 ; 
   reg __411356_411356;
   reg _411357_411357 ; 
   reg __411357_411357;
   reg _411358_411358 ; 
   reg __411358_411358;
   reg _411359_411359 ; 
   reg __411359_411359;
   reg _411360_411360 ; 
   reg __411360_411360;
   reg _411361_411361 ; 
   reg __411361_411361;
   reg _411362_411362 ; 
   reg __411362_411362;
   reg _411363_411363 ; 
   reg __411363_411363;
   reg _411364_411364 ; 
   reg __411364_411364;
   reg _411365_411365 ; 
   reg __411365_411365;
   reg _411366_411366 ; 
   reg __411366_411366;
   reg _411367_411367 ; 
   reg __411367_411367;
   reg _411368_411368 ; 
   reg __411368_411368;
   reg _411369_411369 ; 
   reg __411369_411369;
   reg _411370_411370 ; 
   reg __411370_411370;
   reg _411371_411371 ; 
   reg __411371_411371;
   reg _411372_411372 ; 
   reg __411372_411372;
   reg _411373_411373 ; 
   reg __411373_411373;
   reg _411374_411374 ; 
   reg __411374_411374;
   reg _411375_411375 ; 
   reg __411375_411375;
   reg _411376_411376 ; 
   reg __411376_411376;
   reg _411377_411377 ; 
   reg __411377_411377;
   reg _411378_411378 ; 
   reg __411378_411378;
   reg _411379_411379 ; 
   reg __411379_411379;
   reg _411380_411380 ; 
   reg __411380_411380;
   reg _411381_411381 ; 
   reg __411381_411381;
   reg _411382_411382 ; 
   reg __411382_411382;
   reg _411383_411383 ; 
   reg __411383_411383;
   reg _411384_411384 ; 
   reg __411384_411384;
   reg _411385_411385 ; 
   reg __411385_411385;
   reg _411386_411386 ; 
   reg __411386_411386;
   reg _411387_411387 ; 
   reg __411387_411387;
   reg _411388_411388 ; 
   reg __411388_411388;
   reg _411389_411389 ; 
   reg __411389_411389;
   reg _411390_411390 ; 
   reg __411390_411390;
   reg _411391_411391 ; 
   reg __411391_411391;
   reg _411392_411392 ; 
   reg __411392_411392;
   reg _411393_411393 ; 
   reg __411393_411393;
   reg _411394_411394 ; 
   reg __411394_411394;
   reg _411395_411395 ; 
   reg __411395_411395;
   reg _411396_411396 ; 
   reg __411396_411396;
   reg _411397_411397 ; 
   reg __411397_411397;
   reg _411398_411398 ; 
   reg __411398_411398;
   reg _411399_411399 ; 
   reg __411399_411399;
   reg _411400_411400 ; 
   reg __411400_411400;
   reg _411401_411401 ; 
   reg __411401_411401;
   reg _411402_411402 ; 
   reg __411402_411402;
   reg _411403_411403 ; 
   reg __411403_411403;
   reg _411404_411404 ; 
   reg __411404_411404;
   reg _411405_411405 ; 
   reg __411405_411405;
   reg _411406_411406 ; 
   reg __411406_411406;
   reg _411407_411407 ; 
   reg __411407_411407;
   reg _411408_411408 ; 
   reg __411408_411408;
   reg _411409_411409 ; 
   reg __411409_411409;
   reg _411410_411410 ; 
   reg __411410_411410;
   reg _411411_411411 ; 
   reg __411411_411411;
   reg _411412_411412 ; 
   reg __411412_411412;
   reg _411413_411413 ; 
   reg __411413_411413;
   reg _411414_411414 ; 
   reg __411414_411414;
   reg _411415_411415 ; 
   reg __411415_411415;
   reg _411416_411416 ; 
   reg __411416_411416;
   reg _411417_411417 ; 
   reg __411417_411417;
   reg _411418_411418 ; 
   reg __411418_411418;
   reg _411419_411419 ; 
   reg __411419_411419;
   reg _411420_411420 ; 
   reg __411420_411420;
   reg _411421_411421 ; 
   reg __411421_411421;
   reg _411422_411422 ; 
   reg __411422_411422;
   reg _411423_411423 ; 
   reg __411423_411423;
   reg _411424_411424 ; 
   reg __411424_411424;
   reg _411425_411425 ; 
   reg __411425_411425;
   reg _411426_411426 ; 
   reg __411426_411426;
   reg _411427_411427 ; 
   reg __411427_411427;
   reg _411428_411428 ; 
   reg __411428_411428;
   reg _411429_411429 ; 
   reg __411429_411429;
   reg _411430_411430 ; 
   reg __411430_411430;
   reg _411431_411431 ; 
   reg __411431_411431;
   reg _411432_411432 ; 
   reg __411432_411432;
   reg _411433_411433 ; 
   reg __411433_411433;
   reg _411434_411434 ; 
   reg __411434_411434;
   reg _411435_411435 ; 
   reg __411435_411435;
   reg _411436_411436 ; 
   reg __411436_411436;
   reg _411437_411437 ; 
   reg __411437_411437;
   reg _411438_411438 ; 
   reg __411438_411438;
   reg _411439_411439 ; 
   reg __411439_411439;
   reg _411440_411440 ; 
   reg __411440_411440;
   reg _411441_411441 ; 
   reg __411441_411441;
   reg _411442_411442 ; 
   reg __411442_411442;
   reg _411443_411443 ; 
   reg __411443_411443;
   reg _411444_411444 ; 
   reg __411444_411444;
   reg _411445_411445 ; 
   reg __411445_411445;
   reg _411446_411446 ; 
   reg __411446_411446;
   reg _411447_411447 ; 
   reg __411447_411447;
   reg _411448_411448 ; 
   reg __411448_411448;
   reg _411449_411449 ; 
   reg __411449_411449;
   reg _411450_411450 ; 
   reg __411450_411450;
   reg _411451_411451 ; 
   reg __411451_411451;
   reg _411452_411452 ; 
   reg __411452_411452;
   reg _411453_411453 ; 
   reg __411453_411453;
   reg _411454_411454 ; 
   reg __411454_411454;
   reg _411455_411455 ; 
   reg __411455_411455;
   reg _411456_411456 ; 
   reg __411456_411456;
   reg _411457_411457 ; 
   reg __411457_411457;
   reg _411458_411458 ; 
   reg __411458_411458;
   reg _411459_411459 ; 
   reg __411459_411459;
   reg _411460_411460 ; 
   reg __411460_411460;
   reg _411461_411461 ; 
   reg __411461_411461;
   reg _411462_411462 ; 
   reg __411462_411462;
   reg _411463_411463 ; 
   reg __411463_411463;
   reg _411464_411464 ; 
   reg __411464_411464;
   reg _411465_411465 ; 
   reg __411465_411465;
   reg _411466_411466 ; 
   reg __411466_411466;
   reg _411467_411467 ; 
   reg __411467_411467;
   reg _411468_411468 ; 
   reg __411468_411468;
   reg _411469_411469 ; 
   reg __411469_411469;
   reg _411470_411470 ; 
   reg __411470_411470;
   reg _411471_411471 ; 
   reg __411471_411471;
   reg _411472_411472 ; 
   reg __411472_411472;
   reg _411473_411473 ; 
   reg __411473_411473;
   reg _411474_411474 ; 
   reg __411474_411474;
   reg _411475_411475 ; 
   reg __411475_411475;
   reg _411476_411476 ; 
   reg __411476_411476;
   reg _411477_411477 ; 
   reg __411477_411477;
   reg _411478_411478 ; 
   reg __411478_411478;
   reg _411479_411479 ; 
   reg __411479_411479;
   reg _411480_411480 ; 
   reg __411480_411480;
   reg _411481_411481 ; 
   reg __411481_411481;
   reg _411482_411482 ; 
   reg __411482_411482;
   reg _411483_411483 ; 
   reg __411483_411483;
   reg _411484_411484 ; 
   reg __411484_411484;
   reg _411485_411485 ; 
   reg __411485_411485;
   reg _411486_411486 ; 
   reg __411486_411486;
   reg _411487_411487 ; 
   reg __411487_411487;
   reg _411488_411488 ; 
   reg __411488_411488;
   reg _411489_411489 ; 
   reg __411489_411489;
   reg _411490_411490 ; 
   reg __411490_411490;
   reg _411491_411491 ; 
   reg __411491_411491;
   reg _411492_411492 ; 
   reg __411492_411492;
   reg _411493_411493 ; 
   reg __411493_411493;
   reg _411494_411494 ; 
   reg __411494_411494;
   reg _411495_411495 ; 
   reg __411495_411495;
   reg _411496_411496 ; 
   reg __411496_411496;
   reg _411497_411497 ; 
   reg __411497_411497;
   reg _411498_411498 ; 
   reg __411498_411498;
   reg _411499_411499 ; 
   reg __411499_411499;
   reg _411500_411500 ; 
   reg __411500_411500;
   reg _411501_411501 ; 
   reg __411501_411501;
   reg _411502_411502 ; 
   reg __411502_411502;
   reg _411503_411503 ; 
   reg __411503_411503;
   reg _411504_411504 ; 
   reg __411504_411504;
   reg _411505_411505 ; 
   reg __411505_411505;
   reg _411506_411506 ; 
   reg __411506_411506;
   reg _411507_411507 ; 
   reg __411507_411507;
   reg _411508_411508 ; 
   reg __411508_411508;
   reg _411509_411509 ; 
   reg __411509_411509;
   reg _411510_411510 ; 
   reg __411510_411510;
   reg _411511_411511 ; 
   reg __411511_411511;
   reg _411512_411512 ; 
   reg __411512_411512;
   reg _411513_411513 ; 
   reg __411513_411513;
   reg _411514_411514 ; 
   reg __411514_411514;
   reg _411515_411515 ; 
   reg __411515_411515;
   reg _411516_411516 ; 
   reg __411516_411516;
   reg _411517_411517 ; 
   reg __411517_411517;
   reg _411518_411518 ; 
   reg __411518_411518;
   reg _411519_411519 ; 
   reg __411519_411519;
   reg _411520_411520 ; 
   reg __411520_411520;
   reg _411521_411521 ; 
   reg __411521_411521;
   reg _411522_411522 ; 
   reg __411522_411522;
   reg _411523_411523 ; 
   reg __411523_411523;
   reg _411524_411524 ; 
   reg __411524_411524;
   reg _411525_411525 ; 
   reg __411525_411525;
   reg _411526_411526 ; 
   reg __411526_411526;
   reg _411527_411527 ; 
   reg __411527_411527;
   reg _411528_411528 ; 
   reg __411528_411528;
   reg _411529_411529 ; 
   reg __411529_411529;
   reg _411530_411530 ; 
   reg __411530_411530;
   reg _411531_411531 ; 
   reg __411531_411531;
   reg _411532_411532 ; 
   reg __411532_411532;
   reg _411533_411533 ; 
   reg __411533_411533;
   reg _411534_411534 ; 
   reg __411534_411534;
   reg _411535_411535 ; 
   reg __411535_411535;
   reg _411536_411536 ; 
   reg __411536_411536;
   reg _411537_411537 ; 
   reg __411537_411537;
   reg _411538_411538 ; 
   reg __411538_411538;
   reg _411539_411539 ; 
   reg __411539_411539;
   reg _411540_411540 ; 
   reg __411540_411540;
   reg _411541_411541 ; 
   reg __411541_411541;
   reg _411542_411542 ; 
   reg __411542_411542;
   reg _411543_411543 ; 
   reg __411543_411543;
   reg _411544_411544 ; 
   reg __411544_411544;
   reg _411545_411545 ; 
   reg __411545_411545;
   reg _411546_411546 ; 
   reg __411546_411546;
   reg _411547_411547 ; 
   reg __411547_411547;
   reg _411548_411548 ; 
   reg __411548_411548;
   reg _411549_411549 ; 
   reg __411549_411549;
   reg _411550_411550 ; 
   reg __411550_411550;
   reg _411551_411551 ; 
   reg __411551_411551;
   reg _411552_411552 ; 
   reg __411552_411552;
   reg _411553_411553 ; 
   reg __411553_411553;
   reg _411554_411554 ; 
   reg __411554_411554;
   reg _411555_411555 ; 
   reg __411555_411555;
   reg _411556_411556 ; 
   reg __411556_411556;
   reg _411557_411557 ; 
   reg __411557_411557;
   reg _411558_411558 ; 
   reg __411558_411558;
   reg _411559_411559 ; 
   reg __411559_411559;
   reg _411560_411560 ; 
   reg __411560_411560;
   reg _411561_411561 ; 
   reg __411561_411561;
   reg _411562_411562 ; 
   reg __411562_411562;
   reg _411563_411563 ; 
   reg __411563_411563;
   reg _411564_411564 ; 
   reg __411564_411564;
   reg _411565_411565 ; 
   reg __411565_411565;
   reg _411566_411566 ; 
   reg __411566_411566;
   reg _411567_411567 ; 
   reg __411567_411567;
   reg _411568_411568 ; 
   reg __411568_411568;
   reg _411569_411569 ; 
   reg __411569_411569;
   reg _411570_411570 ; 
   reg __411570_411570;
   reg _411571_411571 ; 
   reg __411571_411571;
   reg _411572_411572 ; 
   reg __411572_411572;
   reg _411573_411573 ; 
   reg __411573_411573;
   reg _411574_411574 ; 
   reg __411574_411574;
   reg _411575_411575 ; 
   reg __411575_411575;
   reg _411576_411576 ; 
   reg __411576_411576;
   reg _411577_411577 ; 
   reg __411577_411577;
   reg _411578_411578 ; 
   reg __411578_411578;
   reg _411579_411579 ; 
   reg __411579_411579;
   reg _411580_411580 ; 
   reg __411580_411580;
   reg _411581_411581 ; 
   reg __411581_411581;
   reg _411582_411582 ; 
   reg __411582_411582;
   reg _411583_411583 ; 
   reg __411583_411583;
   reg _411584_411584 ; 
   reg __411584_411584;
   reg _411585_411585 ; 
   reg __411585_411585;
   reg _411586_411586 ; 
   reg __411586_411586;
   reg _411587_411587 ; 
   reg __411587_411587;
   reg _411588_411588 ; 
   reg __411588_411588;
   reg _411589_411589 ; 
   reg __411589_411589;
   reg _411590_411590 ; 
   reg __411590_411590;
   reg _411591_411591 ; 
   reg __411591_411591;
   reg _411592_411592 ; 
   reg __411592_411592;
   reg _411593_411593 ; 
   reg __411593_411593;
   reg _411594_411594 ; 
   reg __411594_411594;
   reg _411595_411595 ; 
   reg __411595_411595;
   reg _411596_411596 ; 
   reg __411596_411596;
   reg _411597_411597 ; 
   reg __411597_411597;
   reg _411598_411598 ; 
   reg __411598_411598;
   reg _411599_411599 ; 
   reg __411599_411599;
   reg _411600_411600 ; 
   reg __411600_411600;
   reg _411601_411601 ; 
   reg __411601_411601;
   reg _411602_411602 ; 
   reg __411602_411602;
   reg _411603_411603 ; 
   reg __411603_411603;
   reg _411604_411604 ; 
   reg __411604_411604;
   reg _411605_411605 ; 
   reg __411605_411605;
   reg _411606_411606 ; 
   reg __411606_411606;
   reg _411607_411607 ; 
   reg __411607_411607;
   reg _411608_411608 ; 
   reg __411608_411608;
   reg _411609_411609 ; 
   reg __411609_411609;
   reg _411610_411610 ; 
   reg __411610_411610;
   reg _411611_411611 ; 
   reg __411611_411611;
   reg _411612_411612 ; 
   reg __411612_411612;
   reg _411613_411613 ; 
   reg __411613_411613;
   reg _411614_411614 ; 
   reg __411614_411614;
   reg _411615_411615 ; 
   reg __411615_411615;
   reg _411616_411616 ; 
   reg __411616_411616;
   reg _411617_411617 ; 
   reg __411617_411617;
   reg _411618_411618 ; 
   reg __411618_411618;
   reg _411619_411619 ; 
   reg __411619_411619;
   reg _411620_411620 ; 
   reg __411620_411620;
   reg _411621_411621 ; 
   reg __411621_411621;
   reg _411622_411622 ; 
   reg __411622_411622;
   reg _411623_411623 ; 
   reg __411623_411623;
   reg _411624_411624 ; 
   reg __411624_411624;
   reg _411625_411625 ; 
   reg __411625_411625;
   reg _411626_411626 ; 
   reg __411626_411626;
   reg _411627_411627 ; 
   reg __411627_411627;
   reg _411628_411628 ; 
   reg __411628_411628;
   reg _411629_411629 ; 
   reg __411629_411629;
   reg _411630_411630 ; 
   reg __411630_411630;
   reg _411631_411631 ; 
   reg __411631_411631;
   reg _411632_411632 ; 
   reg __411632_411632;
   reg _411633_411633 ; 
   reg __411633_411633;
   reg _411634_411634 ; 
   reg __411634_411634;
   reg _411635_411635 ; 
   reg __411635_411635;
   reg _411636_411636 ; 
   reg __411636_411636;
   reg _411637_411637 ; 
   reg __411637_411637;
   reg _411638_411638 ; 
   reg __411638_411638;
   reg _411639_411639 ; 
   reg __411639_411639;
   reg _411640_411640 ; 
   reg __411640_411640;
   reg _411641_411641 ; 
   reg __411641_411641;
   reg _411642_411642 ; 
   reg __411642_411642;
   reg _411643_411643 ; 
   reg __411643_411643;
   reg _411644_411644 ; 
   reg __411644_411644;
   reg _411645_411645 ; 
   reg __411645_411645;
   reg _411646_411646 ; 
   reg __411646_411646;
   reg _411647_411647 ; 
   reg __411647_411647;
   reg _411648_411648 ; 
   reg __411648_411648;
   reg _411649_411649 ; 
   reg __411649_411649;
   reg _411650_411650 ; 
   reg __411650_411650;
   reg _411651_411651 ; 
   reg __411651_411651;
   reg _411652_411652 ; 
   reg __411652_411652;
   reg _411653_411653 ; 
   reg __411653_411653;
   reg _411654_411654 ; 
   reg __411654_411654;
   reg _411655_411655 ; 
   reg __411655_411655;
   reg _411656_411656 ; 
   reg __411656_411656;
   reg _411657_411657 ; 
   reg __411657_411657;
   reg _411658_411658 ; 
   reg __411658_411658;
   reg _411659_411659 ; 
   reg __411659_411659;
   reg _411660_411660 ; 
   reg __411660_411660;
   reg _411661_411661 ; 
   reg __411661_411661;
   reg _411662_411662 ; 
   reg __411662_411662;
   reg _411663_411663 ; 
   reg __411663_411663;
   reg _411664_411664 ; 
   reg __411664_411664;
   reg _411665_411665 ; 
   reg __411665_411665;
   reg _411666_411666 ; 
   reg __411666_411666;
   reg _411667_411667 ; 
   reg __411667_411667;
   reg _411668_411668 ; 
   reg __411668_411668;
   reg _411669_411669 ; 
   reg __411669_411669;
   reg _411670_411670 ; 
   reg __411670_411670;
   reg _411671_411671 ; 
   reg __411671_411671;
   reg _411672_411672 ; 
   reg __411672_411672;
   reg _411673_411673 ; 
   reg __411673_411673;
   reg _411674_411674 ; 
   reg __411674_411674;
   reg _411675_411675 ; 
   reg __411675_411675;
   reg _411676_411676 ; 
   reg __411676_411676;
   reg _411677_411677 ; 
   reg __411677_411677;
   reg _411678_411678 ; 
   reg __411678_411678;
   reg _411679_411679 ; 
   reg __411679_411679;
   reg _411680_411680 ; 
   reg __411680_411680;
   reg _411681_411681 ; 
   reg __411681_411681;
   reg _411682_411682 ; 
   reg __411682_411682;
   reg _411683_411683 ; 
   reg __411683_411683;
   reg _411684_411684 ; 
   reg __411684_411684;
   reg _411685_411685 ; 
   reg __411685_411685;
   reg _411686_411686 ; 
   reg __411686_411686;
   reg _411687_411687 ; 
   reg __411687_411687;
   reg _411688_411688 ; 
   reg __411688_411688;
   reg _411689_411689 ; 
   reg __411689_411689;
   reg _411690_411690 ; 
   reg __411690_411690;
   reg _411691_411691 ; 
   reg __411691_411691;
   reg _411692_411692 ; 
   reg __411692_411692;
   reg _411693_411693 ; 
   reg __411693_411693;
   reg _411694_411694 ; 
   reg __411694_411694;
   reg _411695_411695 ; 
   reg __411695_411695;
   reg _411696_411696 ; 
   reg __411696_411696;
   reg _411697_411697 ; 
   reg __411697_411697;
   reg _411698_411698 ; 
   reg __411698_411698;
   reg _411699_411699 ; 
   reg __411699_411699;
   reg _411700_411700 ; 
   reg __411700_411700;
   reg _411701_411701 ; 
   reg __411701_411701;
   reg _411702_411702 ; 
   reg __411702_411702;
   reg _411703_411703 ; 
   reg __411703_411703;
   reg _411704_411704 ; 
   reg __411704_411704;
   reg _411705_411705 ; 
   reg __411705_411705;
   reg _411706_411706 ; 
   reg __411706_411706;
   reg _411707_411707 ; 
   reg __411707_411707;
   reg _411708_411708 ; 
   reg __411708_411708;
   reg _411709_411709 ; 
   reg __411709_411709;
   reg _411710_411710 ; 
   reg __411710_411710;
   reg _411711_411711 ; 
   reg __411711_411711;
   reg _411712_411712 ; 
   reg __411712_411712;
   reg _411713_411713 ; 
   reg __411713_411713;
   reg _411714_411714 ; 
   reg __411714_411714;
   reg _411715_411715 ; 
   reg __411715_411715;
   reg _411716_411716 ; 
   reg __411716_411716;
   reg _411717_411717 ; 
   reg __411717_411717;
   reg _411718_411718 ; 
   reg __411718_411718;
   reg _411719_411719 ; 
   reg __411719_411719;
   reg _411720_411720 ; 
   reg __411720_411720;
   reg _411721_411721 ; 
   reg __411721_411721;
   reg _411722_411722 ; 
   reg __411722_411722;
   reg _411723_411723 ; 
   reg __411723_411723;
   reg _411724_411724 ; 
   reg __411724_411724;
   reg _411725_411725 ; 
   reg __411725_411725;
   reg _411726_411726 ; 
   reg __411726_411726;
   reg _411727_411727 ; 
   reg __411727_411727;
   reg _411728_411728 ; 
   reg __411728_411728;
   reg _411729_411729 ; 
   reg __411729_411729;
   reg _411730_411730 ; 
   reg __411730_411730;
   reg _411731_411731 ; 
   reg __411731_411731;
   reg _411732_411732 ; 
   reg __411732_411732;
   reg _411733_411733 ; 
   reg __411733_411733;
   reg _411734_411734 ; 
   reg __411734_411734;
   reg _411735_411735 ; 
   reg __411735_411735;
   reg _411736_411736 ; 
   reg __411736_411736;
   reg _411737_411737 ; 
   reg __411737_411737;
   reg _411738_411738 ; 
   reg __411738_411738;
   reg _411739_411739 ; 
   reg __411739_411739;
   reg _411740_411740 ; 
   reg __411740_411740;
   reg _411741_411741 ; 
   reg __411741_411741;
   reg _411742_411742 ; 
   reg __411742_411742;
   reg _411743_411743 ; 
   reg __411743_411743;
   reg _411744_411744 ; 
   reg __411744_411744;
   reg _411745_411745 ; 
   reg __411745_411745;
   reg _411746_411746 ; 
   reg __411746_411746;
   reg _411747_411747 ; 
   reg __411747_411747;
   reg _411748_411748 ; 
   reg __411748_411748;
   reg _411749_411749 ; 
   reg __411749_411749;
   reg _411750_411750 ; 
   reg __411750_411750;
   reg _411751_411751 ; 
   reg __411751_411751;
   reg _411752_411752 ; 
   reg __411752_411752;
   reg _411753_411753 ; 
   reg __411753_411753;
   reg _411754_411754 ; 
   reg __411754_411754;
   reg _411755_411755 ; 
   reg __411755_411755;
   reg _411756_411756 ; 
   reg __411756_411756;
   reg _411757_411757 ; 
   reg __411757_411757;
   reg _411758_411758 ; 
   reg __411758_411758;
   reg _411759_411759 ; 
   reg __411759_411759;
   reg _411760_411760 ; 
   reg __411760_411760;
   reg _411761_411761 ; 
   reg __411761_411761;
   reg _411762_411762 ; 
   reg __411762_411762;
   reg _411763_411763 ; 
   reg __411763_411763;
   reg _411764_411764 ; 
   reg __411764_411764;
   reg _411765_411765 ; 
   reg __411765_411765;
   reg _411766_411766 ; 
   reg __411766_411766;
   reg _411767_411767 ; 
   reg __411767_411767;
   reg _411768_411768 ; 
   reg __411768_411768;
   reg _411769_411769 ; 
   reg __411769_411769;
   reg _411770_411770 ; 
   reg __411770_411770;
   reg _411771_411771 ; 
   reg __411771_411771;
   reg _411772_411772 ; 
   reg __411772_411772;
   reg _411773_411773 ; 
   reg __411773_411773;
   reg _411774_411774 ; 
   reg __411774_411774;
   reg _411775_411775 ; 
   reg __411775_411775;
   reg _411776_411776 ; 
   reg __411776_411776;
   reg _411777_411777 ; 
   reg __411777_411777;
   reg _411778_411778 ; 
   reg __411778_411778;
   reg _411779_411779 ; 
   reg __411779_411779;
   reg _411780_411780 ; 
   reg __411780_411780;
   reg _411781_411781 ; 
   reg __411781_411781;
   reg _411782_411782 ; 
   reg __411782_411782;
   reg _411783_411783 ; 
   reg __411783_411783;
   reg _411784_411784 ; 
   reg __411784_411784;
   reg _411785_411785 ; 
   reg __411785_411785;
   reg _411786_411786 ; 
   reg __411786_411786;
   reg _411787_411787 ; 
   reg __411787_411787;
   reg _411788_411788 ; 
   reg __411788_411788;
   reg _411789_411789 ; 
   reg __411789_411789;
   reg _411790_411790 ; 
   reg __411790_411790;
   reg _411791_411791 ; 
   reg __411791_411791;
   reg _411792_411792 ; 
   reg __411792_411792;
   reg _411793_411793 ; 
   reg __411793_411793;
   reg _411794_411794 ; 
   reg __411794_411794;
   reg _411795_411795 ; 
   reg __411795_411795;
   reg _411796_411796 ; 
   reg __411796_411796;
   reg _411797_411797 ; 
   reg __411797_411797;
   reg _411798_411798 ; 
   reg __411798_411798;
   reg _411799_411799 ; 
   reg __411799_411799;
   reg _411800_411800 ; 
   reg __411800_411800;
   reg _411801_411801 ; 
   reg __411801_411801;
   reg _411802_411802 ; 
   reg __411802_411802;
   reg _411803_411803 ; 
   reg __411803_411803;
   reg _411804_411804 ; 
   reg __411804_411804;
   reg _411805_411805 ; 
   reg __411805_411805;
   reg _411806_411806 ; 
   reg __411806_411806;
   reg _411807_411807 ; 
   reg __411807_411807;
   reg _411808_411808 ; 
   reg __411808_411808;
   reg _411809_411809 ; 
   reg __411809_411809;
   reg _411810_411810 ; 
   reg __411810_411810;
   reg _411811_411811 ; 
   reg __411811_411811;
   reg _411812_411812 ; 
   reg __411812_411812;
   reg _411813_411813 ; 
   reg __411813_411813;
   reg _411814_411814 ; 
   reg __411814_411814;
   reg _411815_411815 ; 
   reg __411815_411815;
   reg _411816_411816 ; 
   reg __411816_411816;
   reg _411817_411817 ; 
   reg __411817_411817;
   reg _411818_411818 ; 
   reg __411818_411818;
   reg _411819_411819 ; 
   reg __411819_411819;
   reg _411820_411820 ; 
   reg __411820_411820;
   reg _411821_411821 ; 
   reg __411821_411821;
   reg _411822_411822 ; 
   reg __411822_411822;
   reg _411823_411823 ; 
   reg __411823_411823;
   reg _411824_411824 ; 
   reg __411824_411824;
   reg _411825_411825 ; 
   reg __411825_411825;
   reg _411826_411826 ; 
   reg __411826_411826;
   reg _411827_411827 ; 
   reg __411827_411827;
   reg _411828_411828 ; 
   reg __411828_411828;
   reg _411829_411829 ; 
   reg __411829_411829;
   reg _411830_411830 ; 
   reg __411830_411830;
   reg _411831_411831 ; 
   reg __411831_411831;
   reg _411832_411832 ; 
   reg __411832_411832;
   reg _411833_411833 ; 
   reg __411833_411833;
   reg _411834_411834 ; 
   reg __411834_411834;
   reg _411835_411835 ; 
   reg __411835_411835;
   reg _411836_411836 ; 
   reg __411836_411836;
   reg _411837_411837 ; 
   reg __411837_411837;
   reg _411838_411838 ; 
   reg __411838_411838;
   reg _411839_411839 ; 
   reg __411839_411839;
   reg _411840_411840 ; 
   reg __411840_411840;
   reg _411841_411841 ; 
   reg __411841_411841;
   reg _411842_411842 ; 
   reg __411842_411842;
   reg _411843_411843 ; 
   reg __411843_411843;
   reg _411844_411844 ; 
   reg __411844_411844;
   reg _411845_411845 ; 
   reg __411845_411845;
   reg _411846_411846 ; 
   reg __411846_411846;
   reg _411847_411847 ; 
   reg __411847_411847;
   reg _411848_411848 ; 
   reg __411848_411848;
   reg _411849_411849 ; 
   reg __411849_411849;
   reg _411850_411850 ; 
   reg __411850_411850;
   reg _411851_411851 ; 
   reg __411851_411851;
   reg _411852_411852 ; 
   reg __411852_411852;
   reg _411853_411853 ; 
   reg __411853_411853;
   reg _411854_411854 ; 
   reg __411854_411854;
   reg _411855_411855 ; 
   reg __411855_411855;
   reg _411856_411856 ; 
   reg __411856_411856;
   reg _411857_411857 ; 
   reg __411857_411857;
   reg _411858_411858 ; 
   reg __411858_411858;
   reg _411859_411859 ; 
   reg __411859_411859;
   reg _411860_411860 ; 
   reg __411860_411860;
   reg _411861_411861 ; 
   reg __411861_411861;
   reg _411862_411862 ; 
   reg __411862_411862;
   reg _411863_411863 ; 
   reg __411863_411863;
   reg _411864_411864 ; 
   reg __411864_411864;
   reg _411865_411865 ; 
   reg __411865_411865;
   reg _411866_411866 ; 
   reg __411866_411866;
   reg _411867_411867 ; 
   reg __411867_411867;
   reg _411868_411868 ; 
   reg __411868_411868;
   reg _411869_411869 ; 
   reg __411869_411869;
   reg _411870_411870 ; 
   reg __411870_411870;
   reg _411871_411871 ; 
   reg __411871_411871;
   reg _411872_411872 ; 
   reg __411872_411872;
   reg _411873_411873 ; 
   reg __411873_411873;
   reg _411874_411874 ; 
   reg __411874_411874;
   reg _411875_411875 ; 
   reg __411875_411875;
   reg _411876_411876 ; 
   reg __411876_411876;
   reg _411877_411877 ; 
   reg __411877_411877;
   reg _411878_411878 ; 
   reg __411878_411878;
   reg _411879_411879 ; 
   reg __411879_411879;
   reg _411880_411880 ; 
   reg __411880_411880;
   reg _411881_411881 ; 
   reg __411881_411881;
   reg _411882_411882 ; 
   reg __411882_411882;
   reg _411883_411883 ; 
   reg __411883_411883;
   reg _411884_411884 ; 
   reg __411884_411884;
   reg _411885_411885 ; 
   reg __411885_411885;
   reg _411886_411886 ; 
   reg __411886_411886;
   reg _411887_411887 ; 
   reg __411887_411887;
   reg _411888_411888 ; 
   reg __411888_411888;
   reg _411889_411889 ; 
   reg __411889_411889;
   reg _411890_411890 ; 
   reg __411890_411890;
   reg _411891_411891 ; 
   reg __411891_411891;
   reg _411892_411892 ; 
   reg __411892_411892;
   reg _411893_411893 ; 
   reg __411893_411893;
   reg _411894_411894 ; 
   reg __411894_411894;
   reg _411895_411895 ; 
   reg __411895_411895;
   reg _411896_411896 ; 
   reg __411896_411896;
   reg _411897_411897 ; 
   reg __411897_411897;
   reg _411898_411898 ; 
   reg __411898_411898;
   reg _411899_411899 ; 
   reg __411899_411899;
   reg _411900_411900 ; 
   reg __411900_411900;
   reg _411901_411901 ; 
   reg __411901_411901;
   reg _411902_411902 ; 
   reg __411902_411902;
   reg _411903_411903 ; 
   reg __411903_411903;
   reg _411904_411904 ; 
   reg __411904_411904;
   reg _411905_411905 ; 
   reg __411905_411905;
   reg _411906_411906 ; 
   reg __411906_411906;
   reg _411907_411907 ; 
   reg __411907_411907;
   reg _411908_411908 ; 
   reg __411908_411908;
   reg _411909_411909 ; 
   reg __411909_411909;
   reg _411910_411910 ; 
   reg __411910_411910;
   reg _411911_411911 ; 
   reg __411911_411911;
   reg _411912_411912 ; 
   reg __411912_411912;
   reg _411913_411913 ; 
   reg __411913_411913;
   reg _411914_411914 ; 
   reg __411914_411914;
   reg _411915_411915 ; 
   reg __411915_411915;
   reg _411916_411916 ; 
   reg __411916_411916;
   reg _411917_411917 ; 
   reg __411917_411917;
   reg _411918_411918 ; 
   reg __411918_411918;
   reg _411919_411919 ; 
   reg __411919_411919;
   reg _411920_411920 ; 
   reg __411920_411920;
   reg _411921_411921 ; 
   reg __411921_411921;
   reg _411922_411922 ; 
   reg __411922_411922;
   reg _411923_411923 ; 
   reg __411923_411923;
   reg _411924_411924 ; 
   reg __411924_411924;
   reg _411925_411925 ; 
   reg __411925_411925;
   reg _411926_411926 ; 
   reg __411926_411926;
   reg _411927_411927 ; 
   reg __411927_411927;
   reg _411928_411928 ; 
   reg __411928_411928;
   reg _411929_411929 ; 
   reg __411929_411929;
   reg _411930_411930 ; 
   reg __411930_411930;
   reg _411931_411931 ; 
   reg __411931_411931;
   reg _411932_411932 ; 
   reg __411932_411932;
   reg _411933_411933 ; 
   reg __411933_411933;
   reg _411934_411934 ; 
   reg __411934_411934;
   reg _411935_411935 ; 
   reg __411935_411935;
   reg _411936_411936 ; 
   reg __411936_411936;
   reg _411937_411937 ; 
   reg __411937_411937;
   reg _411938_411938 ; 
   reg __411938_411938;
   reg _411939_411939 ; 
   reg __411939_411939;
   reg _411940_411940 ; 
   reg __411940_411940;
   reg _411941_411941 ; 
   reg __411941_411941;
   reg _411942_411942 ; 
   reg __411942_411942;
   reg _411943_411943 ; 
   reg __411943_411943;
   reg _411944_411944 ; 
   reg __411944_411944;
   reg _411945_411945 ; 
   reg __411945_411945;
   reg _411946_411946 ; 
   reg __411946_411946;
   reg _411947_411947 ; 
   reg __411947_411947;
   reg _411948_411948 ; 
   reg __411948_411948;
   reg _411949_411949 ; 
   reg __411949_411949;
   reg _411950_411950 ; 
   reg __411950_411950;
   reg _411951_411951 ; 
   reg __411951_411951;
   reg _411952_411952 ; 
   reg __411952_411952;
   reg _411953_411953 ; 
   reg __411953_411953;
   reg _411954_411954 ; 
   reg __411954_411954;
   reg _411955_411955 ; 
   reg __411955_411955;
   reg _411956_411956 ; 
   reg __411956_411956;
   reg _411957_411957 ; 
   reg __411957_411957;
   reg _411958_411958 ; 
   reg __411958_411958;
   reg _411959_411959 ; 
   reg __411959_411959;
   reg _411960_411960 ; 
   reg __411960_411960;
   reg _411961_411961 ; 
   reg __411961_411961;
   reg _411962_411962 ; 
   reg __411962_411962;
   reg _411963_411963 ; 
   reg __411963_411963;
   reg _411964_411964 ; 
   reg __411964_411964;
   reg _411965_411965 ; 
   reg __411965_411965;
   reg _411966_411966 ; 
   reg __411966_411966;
   reg _411967_411967 ; 
   reg __411967_411967;
   reg _411968_411968 ; 
   reg __411968_411968;
   reg _411969_411969 ; 
   reg __411969_411969;
   reg _411970_411970 ; 
   reg __411970_411970;
   reg _411971_411971 ; 
   reg __411971_411971;
   reg _411972_411972 ; 
   reg __411972_411972;
   reg _411973_411973 ; 
   reg __411973_411973;
   reg _411974_411974 ; 
   reg __411974_411974;
   reg _411975_411975 ; 
   reg __411975_411975;
   reg _411976_411976 ; 
   reg __411976_411976;
   reg _411977_411977 ; 
   reg __411977_411977;
   reg _411978_411978 ; 
   reg __411978_411978;
   reg _411979_411979 ; 
   reg __411979_411979;
   reg _411980_411980 ; 
   reg __411980_411980;
   reg _411981_411981 ; 
   reg __411981_411981;
   reg _411982_411982 ; 
   reg __411982_411982;
   reg _411983_411983 ; 
   reg __411983_411983;
   reg _411984_411984 ; 
   reg __411984_411984;
   reg _411985_411985 ; 
   reg __411985_411985;
   reg _411986_411986 ; 
   reg __411986_411986;
   reg _411987_411987 ; 
   reg __411987_411987;
   reg _411988_411988 ; 
   reg __411988_411988;
   reg _411989_411989 ; 
   reg __411989_411989;
   reg _411990_411990 ; 
   reg __411990_411990;
   reg _411991_411991 ; 
   reg __411991_411991;
   reg _411992_411992 ; 
   reg __411992_411992;
   reg _411993_411993 ; 
   reg __411993_411993;
   reg _411994_411994 ; 
   reg __411994_411994;
   reg _411995_411995 ; 
   reg __411995_411995;
   reg _411996_411996 ; 
   reg __411996_411996;
   reg _411997_411997 ; 
   reg __411997_411997;
   reg _411998_411998 ; 
   reg __411998_411998;
   reg _411999_411999 ; 
   reg __411999_411999;
   reg _412000_412000 ; 
   reg __412000_412000;
   reg _412001_412001 ; 
   reg __412001_412001;
   reg _412002_412002 ; 
   reg __412002_412002;
   reg _412003_412003 ; 
   reg __412003_412003;
   reg _412004_412004 ; 
   reg __412004_412004;
   reg _412005_412005 ; 
   reg __412005_412005;
   reg _412006_412006 ; 
   reg __412006_412006;
   reg _412007_412007 ; 
   reg __412007_412007;
   reg _412008_412008 ; 
   reg __412008_412008;
   reg _412009_412009 ; 
   reg __412009_412009;
   reg _412010_412010 ; 
   reg __412010_412010;
   reg _412011_412011 ; 
   reg __412011_412011;
   reg _412012_412012 ; 
   reg __412012_412012;
   reg _412013_412013 ; 
   reg __412013_412013;
   reg _412014_412014 ; 
   reg __412014_412014;
   reg _412015_412015 ; 
   reg __412015_412015;
   reg _412016_412016 ; 
   reg __412016_412016;
   reg _412017_412017 ; 
   reg __412017_412017;
   reg _412018_412018 ; 
   reg __412018_412018;
   reg _412019_412019 ; 
   reg __412019_412019;
   reg _412020_412020 ; 
   reg __412020_412020;
   reg _412021_412021 ; 
   reg __412021_412021;
   reg _412022_412022 ; 
   reg __412022_412022;
   reg _412023_412023 ; 
   reg __412023_412023;
   reg _412024_412024 ; 
   reg __412024_412024;
   reg _412025_412025 ; 
   reg __412025_412025;
   reg _412026_412026 ; 
   reg __412026_412026;
   reg _412027_412027 ; 
   reg __412027_412027;
   reg _412028_412028 ; 
   reg __412028_412028;
   reg _412029_412029 ; 
   reg __412029_412029;
   reg _412030_412030 ; 
   reg __412030_412030;
   reg _412031_412031 ; 
   reg __412031_412031;
   reg _412032_412032 ; 
   reg __412032_412032;
   reg _412033_412033 ; 
   reg __412033_412033;
   reg _412034_412034 ; 
   reg __412034_412034;
   reg _412035_412035 ; 
   reg __412035_412035;
   reg _412036_412036 ; 
   reg __412036_412036;
   reg _412037_412037 ; 
   reg __412037_412037;
   reg _412038_412038 ; 
   reg __412038_412038;
   reg _412039_412039 ; 
   reg __412039_412039;
   reg _412040_412040 ; 
   reg __412040_412040;
   reg _412041_412041 ; 
   reg __412041_412041;
   reg _412042_412042 ; 
   reg __412042_412042;
   reg _412043_412043 ; 
   reg __412043_412043;
   reg _412044_412044 ; 
   reg __412044_412044;
   reg _412045_412045 ; 
   reg __412045_412045;
   reg _412046_412046 ; 
   reg __412046_412046;
   reg _412047_412047 ; 
   reg __412047_412047;
   reg _412048_412048 ; 
   reg __412048_412048;
   reg _412049_412049 ; 
   reg __412049_412049;
   reg _412050_412050 ; 
   reg __412050_412050;
   reg _412051_412051 ; 
   reg __412051_412051;
   reg _412052_412052 ; 
   reg __412052_412052;
   reg _412053_412053 ; 
   reg __412053_412053;
   reg _412054_412054 ; 
   reg __412054_412054;
   reg _412055_412055 ; 
   reg __412055_412055;
   reg _412056_412056 ; 
   reg __412056_412056;
   reg _412057_412057 ; 
   reg __412057_412057;
   reg _412058_412058 ; 
   reg __412058_412058;
   reg _412059_412059 ; 
   reg __412059_412059;
   reg _412060_412060 ; 
   reg __412060_412060;
   reg _412061_412061 ; 
   reg __412061_412061;
   reg _412062_412062 ; 
   reg __412062_412062;
   reg _412063_412063 ; 
   reg __412063_412063;
   reg _412064_412064 ; 
   reg __412064_412064;
   reg _412065_412065 ; 
   reg __412065_412065;
   reg _412066_412066 ; 
   reg __412066_412066;
   reg _412067_412067 ; 
   reg __412067_412067;
   reg _412068_412068 ; 
   reg __412068_412068;
   reg _412069_412069 ; 
   reg __412069_412069;
   reg _412070_412070 ; 
   reg __412070_412070;
   reg _412071_412071 ; 
   reg __412071_412071;
   reg _412072_412072 ; 
   reg __412072_412072;
   reg _412073_412073 ; 
   reg __412073_412073;
   reg _412074_412074 ; 
   reg __412074_412074;
   reg _412075_412075 ; 
   reg __412075_412075;
   reg _412076_412076 ; 
   reg __412076_412076;
   reg _412077_412077 ; 
   reg __412077_412077;
   reg _412078_412078 ; 
   reg __412078_412078;
   reg _412079_412079 ; 
   reg __412079_412079;
   reg _412080_412080 ; 
   reg __412080_412080;
   reg _412081_412081 ; 
   reg __412081_412081;
   reg _412082_412082 ; 
   reg __412082_412082;
   reg _412083_412083 ; 
   reg __412083_412083;
   reg _412084_412084 ; 
   reg __412084_412084;
   reg _412085_412085 ; 
   reg __412085_412085;
   reg _412086_412086 ; 
   reg __412086_412086;
   reg _412087_412087 ; 
   reg __412087_412087;
   reg _412088_412088 ; 
   reg __412088_412088;
   reg _412089_412089 ; 
   reg __412089_412089;
   reg _412090_412090 ; 
   reg __412090_412090;
   reg _412091_412091 ; 
   reg __412091_412091;
   reg _412092_412092 ; 
   reg __412092_412092;
   reg _412093_412093 ; 
   reg __412093_412093;
   reg _412094_412094 ; 
   reg __412094_412094;
   reg _412095_412095 ; 
   reg __412095_412095;
   reg _412096_412096 ; 
   reg __412096_412096;
   reg _412097_412097 ; 
   reg __412097_412097;
   reg _412098_412098 ; 
   reg __412098_412098;
   reg _412099_412099 ; 
   reg __412099_412099;
   reg _412100_412100 ; 
   reg __412100_412100;
   reg _412101_412101 ; 
   reg __412101_412101;
   reg _412102_412102 ; 
   reg __412102_412102;
   reg _412103_412103 ; 
   reg __412103_412103;
   reg _412104_412104 ; 
   reg __412104_412104;
   reg _412105_412105 ; 
   reg __412105_412105;
   reg _412106_412106 ; 
   reg __412106_412106;
   reg _412107_412107 ; 
   reg __412107_412107;
   reg _412108_412108 ; 
   reg __412108_412108;
   reg _412109_412109 ; 
   reg __412109_412109;
   reg _412110_412110 ; 
   reg __412110_412110;
   reg _412111_412111 ; 
   reg __412111_412111;
   reg _412112_412112 ; 
   reg __412112_412112;
   reg _412113_412113 ; 
   reg __412113_412113;
   reg _412114_412114 ; 
   reg __412114_412114;
   reg _412115_412115 ; 
   reg __412115_412115;
   reg _412116_412116 ; 
   reg __412116_412116;
   reg _412117_412117 ; 
   reg __412117_412117;
   reg _412118_412118 ; 
   reg __412118_412118;
   reg _412119_412119 ; 
   reg __412119_412119;
   reg _412120_412120 ; 
   reg __412120_412120;
   reg _412121_412121 ; 
   reg __412121_412121;
   reg _412122_412122 ; 
   reg __412122_412122;
   reg _412123_412123 ; 
   reg __412123_412123;
   reg _412124_412124 ; 
   reg __412124_412124;
   reg _412125_412125 ; 
   reg __412125_412125;
   reg _412126_412126 ; 
   reg __412126_412126;
   reg _412127_412127 ; 
   reg __412127_412127;
   reg _412128_412128 ; 
   reg __412128_412128;
   reg _412129_412129 ; 
   reg __412129_412129;
   reg _412130_412130 ; 
   reg __412130_412130;
   reg _412131_412131 ; 
   reg __412131_412131;
   reg _412132_412132 ; 
   reg __412132_412132;
   reg _412133_412133 ; 
   reg __412133_412133;
   reg _412134_412134 ; 
   reg __412134_412134;
   reg _412135_412135 ; 
   reg __412135_412135;
   reg _412136_412136 ; 
   reg __412136_412136;
   reg _412137_412137 ; 
   reg __412137_412137;
   reg _412138_412138 ; 
   reg __412138_412138;
   reg _412139_412139 ; 
   reg __412139_412139;
   reg _412140_412140 ; 
   reg __412140_412140;
   reg _412141_412141 ; 
   reg __412141_412141;
   reg _412142_412142 ; 
   reg __412142_412142;
   reg _412143_412143 ; 
   reg __412143_412143;
   reg _412144_412144 ; 
   reg __412144_412144;
   reg _412145_412145 ; 
   reg __412145_412145;
   reg _412146_412146 ; 
   reg __412146_412146;
   reg _412147_412147 ; 
   reg __412147_412147;
   reg _412148_412148 ; 
   reg __412148_412148;
   reg _412149_412149 ; 
   reg __412149_412149;
   reg _412150_412150 ; 
   reg __412150_412150;
   reg _412151_412151 ; 
   reg __412151_412151;
   reg _412152_412152 ; 
   reg __412152_412152;
   reg _412153_412153 ; 
   reg __412153_412153;
   reg _412154_412154 ; 
   reg __412154_412154;
   reg _412155_412155 ; 
   reg __412155_412155;
   reg _412156_412156 ; 
   reg __412156_412156;
   reg _412157_412157 ; 
   reg __412157_412157;
   reg _412158_412158 ; 
   reg __412158_412158;
   reg _412159_412159 ; 
   reg __412159_412159;
   reg _412160_412160 ; 
   reg __412160_412160;
   reg _412161_412161 ; 
   reg __412161_412161;
   reg _412162_412162 ; 
   reg __412162_412162;
   reg _412163_412163 ; 
   reg __412163_412163;
   reg _412164_412164 ; 
   reg __412164_412164;
   reg _412165_412165 ; 
   reg __412165_412165;
   reg _412166_412166 ; 
   reg __412166_412166;
   reg _412167_412167 ; 
   reg __412167_412167;
   reg _412168_412168 ; 
   reg __412168_412168;
   reg _412169_412169 ; 
   reg __412169_412169;
   reg _412170_412170 ; 
   reg __412170_412170;
   reg _412171_412171 ; 
   reg __412171_412171;
   reg _412172_412172 ; 
   reg __412172_412172;
   reg _412173_412173 ; 
   reg __412173_412173;
   reg _412174_412174 ; 
   reg __412174_412174;
   reg _412175_412175 ; 
   reg __412175_412175;
   reg _412176_412176 ; 
   reg __412176_412176;
   reg _412177_412177 ; 
   reg __412177_412177;
   reg _412178_412178 ; 
   reg __412178_412178;
   reg _412179_412179 ; 
   reg __412179_412179;
   reg _412180_412180 ; 
   reg __412180_412180;
   reg _412181_412181 ; 
   reg __412181_412181;
   reg _412182_412182 ; 
   reg __412182_412182;
   reg _412183_412183 ; 
   reg __412183_412183;
   reg _412184_412184 ; 
   reg __412184_412184;
   reg _412185_412185 ; 
   reg __412185_412185;
   reg _412186_412186 ; 
   reg __412186_412186;
   reg _412187_412187 ; 
   reg __412187_412187;
   reg _412188_412188 ; 
   reg __412188_412188;
   reg _412189_412189 ; 
   reg __412189_412189;
   reg _412190_412190 ; 
   reg __412190_412190;
   reg _412191_412191 ; 
   reg __412191_412191;
   reg _412192_412192 ; 
   reg __412192_412192;
   reg _412193_412193 ; 
   reg __412193_412193;
   reg _412194_412194 ; 
   reg __412194_412194;
   reg _412195_412195 ; 
   reg __412195_412195;
   reg _412196_412196 ; 
   reg __412196_412196;
   reg _412197_412197 ; 
   reg __412197_412197;
   reg _412198_412198 ; 
   reg __412198_412198;
   reg _412199_412199 ; 
   reg __412199_412199;
   reg _412200_412200 ; 
   reg __412200_412200;
   reg _412201_412201 ; 
   reg __412201_412201;
   reg _412202_412202 ; 
   reg __412202_412202;
   reg _412203_412203 ; 
   reg __412203_412203;
   reg _412204_412204 ; 
   reg __412204_412204;
   reg _412205_412205 ; 
   reg __412205_412205;
   reg _412206_412206 ; 
   reg __412206_412206;
   reg _412207_412207 ; 
   reg __412207_412207;
   reg _412208_412208 ; 
   reg __412208_412208;
   reg _412209_412209 ; 
   reg __412209_412209;
   reg _412210_412210 ; 
   reg __412210_412210;
   reg _412211_412211 ; 
   reg __412211_412211;
   reg _412212_412212 ; 
   reg __412212_412212;
   reg _412213_412213 ; 
   reg __412213_412213;
   reg _412214_412214 ; 
   reg __412214_412214;
   reg _412215_412215 ; 
   reg __412215_412215;
   reg _412216_412216 ; 
   reg __412216_412216;
   reg _412217_412217 ; 
   reg __412217_412217;
   reg _412218_412218 ; 
   reg __412218_412218;
   reg _412219_412219 ; 
   reg __412219_412219;
   reg _412220_412220 ; 
   reg __412220_412220;
   reg _412221_412221 ; 
   reg __412221_412221;
   reg _412222_412222 ; 
   reg __412222_412222;
   reg _412223_412223 ; 
   reg __412223_412223;
   reg _412224_412224 ; 
   reg __412224_412224;
   reg _412225_412225 ; 
   reg __412225_412225;
   reg _412226_412226 ; 
   reg __412226_412226;
   reg _412227_412227 ; 
   reg __412227_412227;
   reg _412228_412228 ; 
   reg __412228_412228;
   reg _412229_412229 ; 
   reg __412229_412229;
   reg _412230_412230 ; 
   reg __412230_412230;
   reg _412231_412231 ; 
   reg __412231_412231;
   reg _412232_412232 ; 
   reg __412232_412232;
   reg _412233_412233 ; 
   reg __412233_412233;
   reg _412234_412234 ; 
   reg __412234_412234;
   reg _412235_412235 ; 
   reg __412235_412235;
   reg _412236_412236 ; 
   reg __412236_412236;
   reg _412237_412237 ; 
   reg __412237_412237;
   reg _412238_412238 ; 
   reg __412238_412238;
   reg _412239_412239 ; 
   reg __412239_412239;
   reg _412240_412240 ; 
   reg __412240_412240;
   reg _412241_412241 ; 
   reg __412241_412241;
   reg _412242_412242 ; 
   reg __412242_412242;
   reg _412243_412243 ; 
   reg __412243_412243;
   reg _412244_412244 ; 
   reg __412244_412244;
   reg _412245_412245 ; 
   reg __412245_412245;
   reg _412246_412246 ; 
   reg __412246_412246;
   reg _412247_412247 ; 
   reg __412247_412247;
   reg _412248_412248 ; 
   reg __412248_412248;
   reg _412249_412249 ; 
   reg __412249_412249;
   reg _412250_412250 ; 
   reg __412250_412250;
   reg _412251_412251 ; 
   reg __412251_412251;
   reg _412252_412252 ; 
   reg __412252_412252;
   reg _412253_412253 ; 
   reg __412253_412253;
   reg _412254_412254 ; 
   reg __412254_412254;
   reg _412255_412255 ; 
   reg __412255_412255;
   reg _412256_412256 ; 
   reg __412256_412256;
   reg _412257_412257 ; 
   reg __412257_412257;
   reg _412258_412258 ; 
   reg __412258_412258;
   reg _412259_412259 ; 
   reg __412259_412259;
   reg _412260_412260 ; 
   reg __412260_412260;
   reg _412261_412261 ; 
   reg __412261_412261;
   reg _412262_412262 ; 
   reg __412262_412262;
   reg _412263_412263 ; 
   reg __412263_412263;
   reg _412264_412264 ; 
   reg __412264_412264;
   reg _412265_412265 ; 
   reg __412265_412265;
   reg _412266_412266 ; 
   reg __412266_412266;
   reg _412267_412267 ; 
   reg __412267_412267;
   reg _412268_412268 ; 
   reg __412268_412268;
   reg _412269_412269 ; 
   reg __412269_412269;
   reg _412270_412270 ; 
   reg __412270_412270;
   reg _412271_412271 ; 
   reg __412271_412271;
   reg _412272_412272 ; 
   reg __412272_412272;
   reg _412273_412273 ; 
   reg __412273_412273;
   reg _412274_412274 ; 
   reg __412274_412274;
   reg _412275_412275 ; 
   reg __412275_412275;
   reg _412276_412276 ; 
   reg __412276_412276;
   reg _412277_412277 ; 
   reg __412277_412277;
   reg _412278_412278 ; 
   reg __412278_412278;
   reg _412279_412279 ; 
   reg __412279_412279;
   reg _412280_412280 ; 
   reg __412280_412280;
   reg _412281_412281 ; 
   reg __412281_412281;
   reg _412282_412282 ; 
   reg __412282_412282;
   reg _412283_412283 ; 
   reg __412283_412283;
   reg _412284_412284 ; 
   reg __412284_412284;
   reg _412285_412285 ; 
   reg __412285_412285;
   reg _412286_412286 ; 
   reg __412286_412286;
   reg _412287_412287 ; 
   reg __412287_412287;
   reg _412288_412288 ; 
   reg __412288_412288;
   reg _412289_412289 ; 
   reg __412289_412289;
   reg _412290_412290 ; 
   reg __412290_412290;
   reg _412291_412291 ; 
   reg __412291_412291;
   reg _412292_412292 ; 
   reg __412292_412292;
   reg _412293_412293 ; 
   reg __412293_412293;
   reg _412294_412294 ; 
   reg __412294_412294;
   reg _412295_412295 ; 
   reg __412295_412295;
   reg _412296_412296 ; 
   reg __412296_412296;
   reg _412297_412297 ; 
   reg __412297_412297;
   reg _412298_412298 ; 
   reg __412298_412298;
   reg _412299_412299 ; 
   reg __412299_412299;
   reg _412300_412300 ; 
   reg __412300_412300;
   reg _412301_412301 ; 
   reg __412301_412301;
   reg _412302_412302 ; 
   reg __412302_412302;
   reg _412303_412303 ; 
   reg __412303_412303;
   reg _412304_412304 ; 
   reg __412304_412304;
   reg _412305_412305 ; 
   reg __412305_412305;
   reg _412306_412306 ; 
   reg __412306_412306;
   reg _412307_412307 ; 
   reg __412307_412307;
   reg _412308_412308 ; 
   reg __412308_412308;
   reg _412309_412309 ; 
   reg __412309_412309;
   reg _412310_412310 ; 
   reg __412310_412310;
   reg _412311_412311 ; 
   reg __412311_412311;
   reg _412312_412312 ; 
   reg __412312_412312;
   reg _412313_412313 ; 
   reg __412313_412313;
   reg _412314_412314 ; 
   reg __412314_412314;
   reg _412315_412315 ; 
   reg __412315_412315;
   reg _412316_412316 ; 
   reg __412316_412316;
   reg _412317_412317 ; 
   reg __412317_412317;
   reg _412318_412318 ; 
   reg __412318_412318;
   reg _412319_412319 ; 
   reg __412319_412319;
   reg _412320_412320 ; 
   reg __412320_412320;
   reg _412321_412321 ; 
   reg __412321_412321;
   reg _412322_412322 ; 
   reg __412322_412322;
   reg _412323_412323 ; 
   reg __412323_412323;
   reg _412324_412324 ; 
   reg __412324_412324;
   reg _412325_412325 ; 
   reg __412325_412325;
   reg _412326_412326 ; 
   reg __412326_412326;
   reg _412327_412327 ; 
   reg __412327_412327;
   reg _412328_412328 ; 
   reg __412328_412328;
   reg _412329_412329 ; 
   reg __412329_412329;
   reg _412330_412330 ; 
   reg __412330_412330;
   reg _412331_412331 ; 
   reg __412331_412331;
   reg _412332_412332 ; 
   reg __412332_412332;
   reg _412333_412333 ; 
   reg __412333_412333;
   reg _412334_412334 ; 
   reg __412334_412334;
   reg _412335_412335 ; 
   reg __412335_412335;
   reg _412336_412336 ; 
   reg __412336_412336;
   reg _412337_412337 ; 
   reg __412337_412337;
   reg _412338_412338 ; 
   reg __412338_412338;
   reg _412339_412339 ; 
   reg __412339_412339;
   reg _412340_412340 ; 
   reg __412340_412340;
   reg _412341_412341 ; 
   reg __412341_412341;
   reg _412342_412342 ; 
   reg __412342_412342;
   reg _412343_412343 ; 
   reg __412343_412343;
   reg _412344_412344 ; 
   reg __412344_412344;
   reg _412345_412345 ; 
   reg __412345_412345;
   reg _412346_412346 ; 
   reg __412346_412346;
   reg _412347_412347 ; 
   reg __412347_412347;
   reg _412348_412348 ; 
   reg __412348_412348;
   reg _412349_412349 ; 
   reg __412349_412349;
   reg _412350_412350 ; 
   reg __412350_412350;
   reg _412351_412351 ; 
   reg __412351_412351;
   reg _412352_412352 ; 
   reg __412352_412352;
   reg _412353_412353 ; 
   reg __412353_412353;
   reg _412354_412354 ; 
   reg __412354_412354;
   reg _412355_412355 ; 
   reg __412355_412355;
   reg _412356_412356 ; 
   reg __412356_412356;
   reg _412357_412357 ; 
   reg __412357_412357;
   reg _412358_412358 ; 
   reg __412358_412358;
   reg _412359_412359 ; 
   reg __412359_412359;
   reg _412360_412360 ; 
   reg __412360_412360;
   reg _412361_412361 ; 
   reg __412361_412361;
   reg _412362_412362 ; 
   reg __412362_412362;
   reg _412363_412363 ; 
   reg __412363_412363;
   reg _412364_412364 ; 
   reg __412364_412364;
   reg _412365_412365 ; 
   reg __412365_412365;
   reg _412366_412366 ; 
   reg __412366_412366;
   reg _412367_412367 ; 
   reg __412367_412367;
   reg _412368_412368 ; 
   reg __412368_412368;
   reg _412369_412369 ; 
   reg __412369_412369;
   reg _412370_412370 ; 
   reg __412370_412370;
   reg _412371_412371 ; 
   reg __412371_412371;
   reg _412372_412372 ; 
   reg __412372_412372;
   reg _412373_412373 ; 
   reg __412373_412373;
   reg _412374_412374 ; 
   reg __412374_412374;
   reg _412375_412375 ; 
   reg __412375_412375;
   reg _412376_412376 ; 
   reg __412376_412376;
   reg _412377_412377 ; 
   reg __412377_412377;
   reg _412378_412378 ; 
   reg __412378_412378;
   reg _412379_412379 ; 
   reg __412379_412379;
   reg _412380_412380 ; 
   reg __412380_412380;
   reg _412381_412381 ; 
   reg __412381_412381;
   reg _412382_412382 ; 
   reg __412382_412382;
   reg _412383_412383 ; 
   reg __412383_412383;
   reg _412384_412384 ; 
   reg __412384_412384;
   reg _412385_412385 ; 
   reg __412385_412385;
   reg _412386_412386 ; 
   reg __412386_412386;
   reg _412387_412387 ; 
   reg __412387_412387;
   reg _412388_412388 ; 
   reg __412388_412388;
   reg _412389_412389 ; 
   reg __412389_412389;
   reg _412390_412390 ; 
   reg __412390_412390;
   reg _412391_412391 ; 
   reg __412391_412391;
   reg _412392_412392 ; 
   reg __412392_412392;
   reg _412393_412393 ; 
   reg __412393_412393;
   reg _412394_412394 ; 
   reg __412394_412394;
   reg _412395_412395 ; 
   reg __412395_412395;
   reg _412396_412396 ; 
   reg __412396_412396;
   reg _412397_412397 ; 
   reg __412397_412397;
   reg _412398_412398 ; 
   reg __412398_412398;
   reg _412399_412399 ; 
   reg __412399_412399;
   reg _412400_412400 ; 
   reg __412400_412400;
   reg _412401_412401 ; 
   reg __412401_412401;
   reg _412402_412402 ; 
   reg __412402_412402;
   reg _412403_412403 ; 
   reg __412403_412403;
   reg _412404_412404 ; 
   reg __412404_412404;
   reg _412405_412405 ; 
   reg __412405_412405;
   reg _412406_412406 ; 
   reg __412406_412406;
   reg _412407_412407 ; 
   reg __412407_412407;
   reg _412408_412408 ; 
   reg __412408_412408;
   reg _412409_412409 ; 
   reg __412409_412409;
   reg _412410_412410 ; 
   reg __412410_412410;
   reg _412411_412411 ; 
   reg __412411_412411;
   reg _412412_412412 ; 
   reg __412412_412412;
   reg _412413_412413 ; 
   reg __412413_412413;
   reg _412414_412414 ; 
   reg __412414_412414;
   reg _412415_412415 ; 
   reg __412415_412415;
   reg _412416_412416 ; 
   reg __412416_412416;
   reg _412417_412417 ; 
   reg __412417_412417;
   reg _412418_412418 ; 
   reg __412418_412418;
   reg _412419_412419 ; 
   reg __412419_412419;
   reg _412420_412420 ; 
   reg __412420_412420;
   reg _412421_412421 ; 
   reg __412421_412421;
   reg _412422_412422 ; 
   reg __412422_412422;
   reg _412423_412423 ; 
   reg __412423_412423;
   reg _412424_412424 ; 
   reg __412424_412424;
   reg _412425_412425 ; 
   reg __412425_412425;
   reg _412426_412426 ; 
   reg __412426_412426;
   reg _412427_412427 ; 
   reg __412427_412427;
   reg _412428_412428 ; 
   reg __412428_412428;
   reg _412429_412429 ; 
   reg __412429_412429;
   reg _412430_412430 ; 
   reg __412430_412430;
   reg _412431_412431 ; 
   reg __412431_412431;
   reg _412432_412432 ; 
   reg __412432_412432;
   reg _412433_412433 ; 
   reg __412433_412433;
   reg _412434_412434 ; 
   reg __412434_412434;
   reg _412435_412435 ; 
   reg __412435_412435;
   reg _412436_412436 ; 
   reg __412436_412436;
   reg _412437_412437 ; 
   reg __412437_412437;
   reg _412438_412438 ; 
   reg __412438_412438;
   reg _412439_412439 ; 
   reg __412439_412439;
   reg _412440_412440 ; 
   reg __412440_412440;
   reg _412441_412441 ; 
   reg __412441_412441;
   reg _412442_412442 ; 
   reg __412442_412442;
   reg _412443_412443 ; 
   reg __412443_412443;
   reg _412444_412444 ; 
   reg __412444_412444;
   reg _412445_412445 ; 
   reg __412445_412445;
   reg _412446_412446 ; 
   reg __412446_412446;
   reg _412447_412447 ; 
   reg __412447_412447;
   reg _412448_412448 ; 
   reg __412448_412448;
   reg _412449_412449 ; 
   reg __412449_412449;
   reg _412450_412450 ; 
   reg __412450_412450;
   reg _412451_412451 ; 
   reg __412451_412451;
   reg _412452_412452 ; 
   reg __412452_412452;
   reg _412453_412453 ; 
   reg __412453_412453;
   reg _412454_412454 ; 
   reg __412454_412454;
   reg _412455_412455 ; 
   reg __412455_412455;
   reg _412456_412456 ; 
   reg __412456_412456;
   reg _412457_412457 ; 
   reg __412457_412457;
   reg _412458_412458 ; 
   reg __412458_412458;
   reg _412459_412459 ; 
   reg __412459_412459;
   reg _412460_412460 ; 
   reg __412460_412460;
   reg _412461_412461 ; 
   reg __412461_412461;
   reg _412462_412462 ; 
   reg __412462_412462;
   reg _412463_412463 ; 
   reg __412463_412463;
   reg _412464_412464 ; 
   reg __412464_412464;
   reg _412465_412465 ; 
   reg __412465_412465;
   reg _412466_412466 ; 
   reg __412466_412466;
   reg _412467_412467 ; 
   reg __412467_412467;
   reg _412468_412468 ; 
   reg __412468_412468;
   reg _412469_412469 ; 
   reg __412469_412469;
   reg _412470_412470 ; 
   reg __412470_412470;
   reg _412471_412471 ; 
   reg __412471_412471;
   reg _412472_412472 ; 
   reg __412472_412472;
   reg _412473_412473 ; 
   reg __412473_412473;
   reg _412474_412474 ; 
   reg __412474_412474;
   reg _412475_412475 ; 
   reg __412475_412475;
   reg _412476_412476 ; 
   reg __412476_412476;
   reg _412477_412477 ; 
   reg __412477_412477;
   reg _412478_412478 ; 
   reg __412478_412478;
   reg _412479_412479 ; 
   reg __412479_412479;
   reg _412480_412480 ; 
   reg __412480_412480;
   reg _412481_412481 ; 
   reg __412481_412481;
   reg _412482_412482 ; 
   reg __412482_412482;
   reg _412483_412483 ; 
   reg __412483_412483;
   reg _412484_412484 ; 
   reg __412484_412484;
   reg _412485_412485 ; 
   reg __412485_412485;
   reg _412486_412486 ; 
   reg __412486_412486;
   reg _412487_412487 ; 
   reg __412487_412487;
   reg _412488_412488 ; 
   reg __412488_412488;
   reg _412489_412489 ; 
   reg __412489_412489;
   reg _412490_412490 ; 
   reg __412490_412490;
   reg _412491_412491 ; 
   reg __412491_412491;
   reg _412492_412492 ; 
   reg __412492_412492;
   reg _412493_412493 ; 
   reg __412493_412493;
   reg _412494_412494 ; 
   reg __412494_412494;
   reg _412495_412495 ; 
   reg __412495_412495;
   reg _412496_412496 ; 
   reg __412496_412496;
   reg _412497_412497 ; 
   reg __412497_412497;
   reg _412498_412498 ; 
   reg __412498_412498;
   reg _412499_412499 ; 
   reg __412499_412499;
   reg _412500_412500 ; 
   reg __412500_412500;
   reg _412501_412501 ; 
   reg __412501_412501;
   reg _412502_412502 ; 
   reg __412502_412502;
   reg _412503_412503 ; 
   reg __412503_412503;
   reg _412504_412504 ; 
   reg __412504_412504;
   reg _412505_412505 ; 
   reg __412505_412505;
   reg _412506_412506 ; 
   reg __412506_412506;
   reg _412507_412507 ; 
   reg __412507_412507;
   reg _412508_412508 ; 
   reg __412508_412508;
   reg _412509_412509 ; 
   reg __412509_412509;
   reg _412510_412510 ; 
   reg __412510_412510;
   reg _412511_412511 ; 
   reg __412511_412511;
   reg _412512_412512 ; 
   reg __412512_412512;
   reg _412513_412513 ; 
   reg __412513_412513;
   reg _412514_412514 ; 
   reg __412514_412514;
   reg _412515_412515 ; 
   reg __412515_412515;
   reg _412516_412516 ; 
   reg __412516_412516;
   reg _412517_412517 ; 
   reg __412517_412517;
   reg _412518_412518 ; 
   reg __412518_412518;
   reg _412519_412519 ; 
   reg __412519_412519;
   reg _412520_412520 ; 
   reg __412520_412520;
   reg _412521_412521 ; 
   reg __412521_412521;
   reg _412522_412522 ; 
   reg __412522_412522;
   reg _412523_412523 ; 
   reg __412523_412523;
   reg _412524_412524 ; 
   reg __412524_412524;
   reg _412525_412525 ; 
   reg __412525_412525;
   reg _412526_412526 ; 
   reg __412526_412526;
   reg _412527_412527 ; 
   reg __412527_412527;
   reg _412528_412528 ; 
   reg __412528_412528;
   reg _412529_412529 ; 
   reg __412529_412529;
   reg _412530_412530 ; 
   reg __412530_412530;
   reg _412531_412531 ; 
   reg __412531_412531;
   reg _412532_412532 ; 
   reg __412532_412532;
   reg _412533_412533 ; 
   reg __412533_412533;
   reg _412534_412534 ; 
   reg __412534_412534;
   reg _412535_412535 ; 
   reg __412535_412535;
   reg _412536_412536 ; 
   reg __412536_412536;
   reg _412537_412537 ; 
   reg __412537_412537;
   reg _412538_412538 ; 
   reg __412538_412538;
   reg _412539_412539 ; 
   reg __412539_412539;
   reg _412540_412540 ; 
   reg __412540_412540;
   reg _412541_412541 ; 
   reg __412541_412541;
   reg _412542_412542 ; 
   reg __412542_412542;
   reg _412543_412543 ; 
   reg __412543_412543;
   reg _412544_412544 ; 
   reg __412544_412544;
   reg _412545_412545 ; 
   reg __412545_412545;
   reg _412546_412546 ; 
   reg __412546_412546;
   reg _412547_412547 ; 
   reg __412547_412547;
   reg _412548_412548 ; 
   reg __412548_412548;
   reg _412549_412549 ; 
   reg __412549_412549;
   reg _412550_412550 ; 
   reg __412550_412550;
   reg _412551_412551 ; 
   reg __412551_412551;
   reg _412552_412552 ; 
   reg __412552_412552;
   reg _412553_412553 ; 
   reg __412553_412553;
   reg _412554_412554 ; 
   reg __412554_412554;
   reg _412555_412555 ; 
   reg __412555_412555;
   reg _412556_412556 ; 
   reg __412556_412556;
   reg _412557_412557 ; 
   reg __412557_412557;
   reg _412558_412558 ; 
   reg __412558_412558;
   reg _412559_412559 ; 
   reg __412559_412559;
   reg _412560_412560 ; 
   reg __412560_412560;
   reg _412561_412561 ; 
   reg __412561_412561;
   reg _412562_412562 ; 
   reg __412562_412562;
   reg _412563_412563 ; 
   reg __412563_412563;
   reg _412564_412564 ; 
   reg __412564_412564;
   reg _412565_412565 ; 
   reg __412565_412565;
   reg _412566_412566 ; 
   reg __412566_412566;
   reg _412567_412567 ; 
   reg __412567_412567;
   reg _412568_412568 ; 
   reg __412568_412568;
   reg _412569_412569 ; 
   reg __412569_412569;
   reg _412570_412570 ; 
   reg __412570_412570;
   reg _412571_412571 ; 
   reg __412571_412571;
   reg _412572_412572 ; 
   reg __412572_412572;
   reg _412573_412573 ; 
   reg __412573_412573;
   reg _412574_412574 ; 
   reg __412574_412574;
   reg _412575_412575 ; 
   reg __412575_412575;
   reg _412576_412576 ; 
   reg __412576_412576;
   reg _412577_412577 ; 
   reg __412577_412577;
   reg _412578_412578 ; 
   reg __412578_412578;
   reg _412579_412579 ; 
   reg __412579_412579;
   reg _412580_412580 ; 
   reg __412580_412580;
   reg _412581_412581 ; 
   reg __412581_412581;
   reg _412582_412582 ; 
   reg __412582_412582;
   reg _412583_412583 ; 
   reg __412583_412583;
   reg _412584_412584 ; 
   reg __412584_412584;
   reg _412585_412585 ; 
   reg __412585_412585;
   reg _412586_412586 ; 
   reg __412586_412586;
   reg _412587_412587 ; 
   reg __412587_412587;
   reg _412588_412588 ; 
   reg __412588_412588;
   reg _412589_412589 ; 
   reg __412589_412589;
   reg _412590_412590 ; 
   reg __412590_412590;
   reg _412591_412591 ; 
   reg __412591_412591;
   reg _412592_412592 ; 
   reg __412592_412592;
   reg _412593_412593 ; 
   reg __412593_412593;
   reg _412594_412594 ; 
   reg __412594_412594;
   reg _412595_412595 ; 
   reg __412595_412595;
   reg _412596_412596 ; 
   reg __412596_412596;
   reg _412597_412597 ; 
   reg __412597_412597;
   reg _412598_412598 ; 
   reg __412598_412598;
   reg _412599_412599 ; 
   reg __412599_412599;
   reg _412600_412600 ; 
   reg __412600_412600;
   reg _412601_412601 ; 
   reg __412601_412601;
   reg _412602_412602 ; 
   reg __412602_412602;
   reg _412603_412603 ; 
   reg __412603_412603;
   reg _412604_412604 ; 
   reg __412604_412604;
   reg _412605_412605 ; 
   reg __412605_412605;
   reg _412606_412606 ; 
   reg __412606_412606;
   reg _412607_412607 ; 
   reg __412607_412607;
   reg _412608_412608 ; 
   reg __412608_412608;
   reg _412609_412609 ; 
   reg __412609_412609;
   reg _412610_412610 ; 
   reg __412610_412610;
   reg _412611_412611 ; 
   reg __412611_412611;
   reg _412612_412612 ; 
   reg __412612_412612;
   reg _412613_412613 ; 
   reg __412613_412613;
   reg _412614_412614 ; 
   reg __412614_412614;
   reg _412615_412615 ; 
   reg __412615_412615;
   reg _412616_412616 ; 
   reg __412616_412616;
   reg _412617_412617 ; 
   reg __412617_412617;
   reg _412618_412618 ; 
   reg __412618_412618;
   reg _412619_412619 ; 
   reg __412619_412619;
   reg _412620_412620 ; 
   reg __412620_412620;
   reg _412621_412621 ; 
   reg __412621_412621;
   reg _412622_412622 ; 
   reg __412622_412622;
   reg _412623_412623 ; 
   reg __412623_412623;
   reg _412624_412624 ; 
   reg __412624_412624;
   reg _412625_412625 ; 
   reg __412625_412625;
   reg _412626_412626 ; 
   reg __412626_412626;
   reg _412627_412627 ; 
   reg __412627_412627;
   reg _412628_412628 ; 
   reg __412628_412628;
   reg _412629_412629 ; 
   reg __412629_412629;
   reg _412630_412630 ; 
   reg __412630_412630;
   reg _412631_412631 ; 
   reg __412631_412631;
   reg _412632_412632 ; 
   reg __412632_412632;
   reg _412633_412633 ; 
   reg __412633_412633;
   reg _412634_412634 ; 
   reg __412634_412634;
   reg _412635_412635 ; 
   reg __412635_412635;
   reg _412636_412636 ; 
   reg __412636_412636;
   reg _412637_412637 ; 
   reg __412637_412637;
   reg _412638_412638 ; 
   reg __412638_412638;
   reg _412639_412639 ; 
   reg __412639_412639;
   reg _412640_412640 ; 
   reg __412640_412640;
   reg _412641_412641 ; 
   reg __412641_412641;
   reg _412642_412642 ; 
   reg __412642_412642;
   reg _412643_412643 ; 
   reg __412643_412643;
   reg _412644_412644 ; 
   reg __412644_412644;
   reg _412645_412645 ; 
   reg __412645_412645;
   reg _412646_412646 ; 
   reg __412646_412646;
   reg _412647_412647 ; 
   reg __412647_412647;
   reg _412648_412648 ; 
   reg __412648_412648;
   reg _412649_412649 ; 
   reg __412649_412649;
   reg _412650_412650 ; 
   reg __412650_412650;
   reg _412651_412651 ; 
   reg __412651_412651;
   reg _412652_412652 ; 
   reg __412652_412652;
   reg _412653_412653 ; 
   reg __412653_412653;
   reg _412654_412654 ; 
   reg __412654_412654;
   reg _412655_412655 ; 
   reg __412655_412655;
   reg _412656_412656 ; 
   reg __412656_412656;
   reg _412657_412657 ; 
   reg __412657_412657;
   reg _412658_412658 ; 
   reg __412658_412658;
   reg _412659_412659 ; 
   reg __412659_412659;
   reg _412660_412660 ; 
   reg __412660_412660;
   reg _412661_412661 ; 
   reg __412661_412661;
   reg _412662_412662 ; 
   reg __412662_412662;
   reg _412663_412663 ; 
   reg __412663_412663;
   reg _412664_412664 ; 
   reg __412664_412664;
   reg _412665_412665 ; 
   reg __412665_412665;
   reg _412666_412666 ; 
   reg __412666_412666;
   reg _412667_412667 ; 
   reg __412667_412667;
   reg _412668_412668 ; 
   reg __412668_412668;
   reg _412669_412669 ; 
   reg __412669_412669;
   reg _412670_412670 ; 
   reg __412670_412670;
   reg _412671_412671 ; 
   reg __412671_412671;
   reg _412672_412672 ; 
   reg __412672_412672;
   reg _412673_412673 ; 
   reg __412673_412673;
   reg _412674_412674 ; 
   reg __412674_412674;
   reg _412675_412675 ; 
   reg __412675_412675;
   reg _412676_412676 ; 
   reg __412676_412676;
   reg _412677_412677 ; 
   reg __412677_412677;
   reg _412678_412678 ; 
   reg __412678_412678;
   reg _412679_412679 ; 
   reg __412679_412679;
   reg _412680_412680 ; 
   reg __412680_412680;
   reg _412681_412681 ; 
   reg __412681_412681;
   reg _412682_412682 ; 
   reg __412682_412682;
   reg _412683_412683 ; 
   reg __412683_412683;
   reg _412684_412684 ; 
   reg __412684_412684;
   reg _412685_412685 ; 
   reg __412685_412685;
   reg _412686_412686 ; 
   reg __412686_412686;
   reg _412687_412687 ; 
   reg __412687_412687;
   reg _412688_412688 ; 
   reg __412688_412688;
   reg _412689_412689 ; 
   reg __412689_412689;
   reg _412690_412690 ; 
   reg __412690_412690;
   reg _412691_412691 ; 
   reg __412691_412691;
   reg _412692_412692 ; 
   reg __412692_412692;
   reg _412693_412693 ; 
   reg __412693_412693;
   reg _412694_412694 ; 
   reg __412694_412694;
   reg _412695_412695 ; 
   reg __412695_412695;
   reg _412696_412696 ; 
   reg __412696_412696;
   reg _412697_412697 ; 
   reg __412697_412697;
   reg _412698_412698 ; 
   reg __412698_412698;
   reg _412699_412699 ; 
   reg __412699_412699;
   reg _412700_412700 ; 
   reg __412700_412700;
   reg _412701_412701 ; 
   reg __412701_412701;
   reg _412702_412702 ; 
   reg __412702_412702;
   reg _412703_412703 ; 
   reg __412703_412703;
   reg _412704_412704 ; 
   reg __412704_412704;
   reg _412705_412705 ; 
   reg __412705_412705;
   reg _412706_412706 ; 
   reg __412706_412706;
   reg _412707_412707 ; 
   reg __412707_412707;
   reg _412708_412708 ; 
   reg __412708_412708;
   reg _412709_412709 ; 
   reg __412709_412709;
   reg _412710_412710 ; 
   reg __412710_412710;
   reg _412711_412711 ; 
   reg __412711_412711;
   reg _412712_412712 ; 
   reg __412712_412712;
   reg _412713_412713 ; 
   reg __412713_412713;
   reg _412714_412714 ; 
   reg __412714_412714;
   reg _412715_412715 ; 
   reg __412715_412715;
   reg _412716_412716 ; 
   reg __412716_412716;
   reg _412717_412717 ; 
   reg __412717_412717;
   reg _412718_412718 ; 
   reg __412718_412718;
   reg _412719_412719 ; 
   reg __412719_412719;
   reg _412720_412720 ; 
   reg __412720_412720;
   reg _412721_412721 ; 
   reg __412721_412721;
   reg _412722_412722 ; 
   reg __412722_412722;
   reg _412723_412723 ; 
   reg __412723_412723;
   reg _412724_412724 ; 
   reg __412724_412724;
   reg _412725_412725 ; 
   reg __412725_412725;
   reg _412726_412726 ; 
   reg __412726_412726;
   reg _412727_412727 ; 
   reg __412727_412727;
   reg _412728_412728 ; 
   reg __412728_412728;
   reg _412729_412729 ; 
   reg __412729_412729;
   reg _412730_412730 ; 
   reg __412730_412730;
   reg _412731_412731 ; 
   reg __412731_412731;
   reg _412732_412732 ; 
   reg __412732_412732;
   reg _412733_412733 ; 
   reg __412733_412733;
   reg _412734_412734 ; 
   reg __412734_412734;
   reg _412735_412735 ; 
   reg __412735_412735;
   reg _412736_412736 ; 
   reg __412736_412736;
   reg _412737_412737 ; 
   reg __412737_412737;
   reg _412738_412738 ; 
   reg __412738_412738;
   reg _412739_412739 ; 
   reg __412739_412739;
   reg _412740_412740 ; 
   reg __412740_412740;
   reg _412741_412741 ; 
   reg __412741_412741;
   reg _412742_412742 ; 
   reg __412742_412742;
   reg _412743_412743 ; 
   reg __412743_412743;
   reg _412744_412744 ; 
   reg __412744_412744;
   reg _412745_412745 ; 
   reg __412745_412745;
   reg _412746_412746 ; 
   reg __412746_412746;
   reg _412747_412747 ; 
   reg __412747_412747;
   reg _412748_412748 ; 
   reg __412748_412748;
   reg _412749_412749 ; 
   reg __412749_412749;
   reg _412750_412750 ; 
   reg __412750_412750;
   reg _412751_412751 ; 
   reg __412751_412751;
   reg _412752_412752 ; 
   reg __412752_412752;
   reg _412753_412753 ; 
   reg __412753_412753;
   reg _412754_412754 ; 
   reg __412754_412754;
   reg _412755_412755 ; 
   reg __412755_412755;
   reg _412756_412756 ; 
   reg __412756_412756;
   reg _412757_412757 ; 
   reg __412757_412757;
   reg _412758_412758 ; 
   reg __412758_412758;
   reg _412759_412759 ; 
   reg __412759_412759;
   reg _412760_412760 ; 
   reg __412760_412760;
   reg _412761_412761 ; 
   reg __412761_412761;
   reg _412762_412762 ; 
   reg __412762_412762;
   reg _412763_412763 ; 
   reg __412763_412763;
   reg _412764_412764 ; 
   reg __412764_412764;
   reg _412765_412765 ; 
   reg __412765_412765;
   reg _412766_412766 ; 
   reg __412766_412766;
   reg _412767_412767 ; 
   reg __412767_412767;
   reg _412768_412768 ; 
   reg __412768_412768;
   reg _412769_412769 ; 
   reg __412769_412769;
   reg _412770_412770 ; 
   reg __412770_412770;
   reg _412771_412771 ; 
   reg __412771_412771;
   reg _412772_412772 ; 
   reg __412772_412772;
   reg _412773_412773 ; 
   reg __412773_412773;
   reg _412774_412774 ; 
   reg __412774_412774;
   reg _412775_412775 ; 
   reg __412775_412775;
   reg _412776_412776 ; 
   reg __412776_412776;
   reg _412777_412777 ; 
   reg __412777_412777;
   reg _412778_412778 ; 
   reg __412778_412778;
   reg _412779_412779 ; 
   reg __412779_412779;
   reg _412780_412780 ; 
   reg __412780_412780;
   reg _412781_412781 ; 
   reg __412781_412781;
   reg _412782_412782 ; 
   reg __412782_412782;
   reg _412783_412783 ; 
   reg __412783_412783;
   reg _412784_412784 ; 
   reg __412784_412784;
   reg _412785_412785 ; 
   reg __412785_412785;
   reg _412786_412786 ; 
   reg __412786_412786;
   reg _412787_412787 ; 
   reg __412787_412787;
   reg _412788_412788 ; 
   reg __412788_412788;
   reg _412789_412789 ; 
   reg __412789_412789;
   reg _412790_412790 ; 
   reg __412790_412790;
   reg _412791_412791 ; 
   reg __412791_412791;
   reg _412792_412792 ; 
   reg __412792_412792;
   reg _412793_412793 ; 
   reg __412793_412793;
   reg _412794_412794 ; 
   reg __412794_412794;
   reg _412795_412795 ; 
   reg __412795_412795;
   reg _412796_412796 ; 
   reg __412796_412796;
   reg _412797_412797 ; 
   reg __412797_412797;
   reg _412798_412798 ; 
   reg __412798_412798;
   reg _412799_412799 ; 
   reg __412799_412799;
   reg _412800_412800 ; 
   reg __412800_412800;
   reg _412801_412801 ; 
   reg __412801_412801;
   reg _412802_412802 ; 
   reg __412802_412802;
   reg _412803_412803 ; 
   reg __412803_412803;
   reg _412804_412804 ; 
   reg __412804_412804;
   reg _412805_412805 ; 
   reg __412805_412805;
   reg _412806_412806 ; 
   reg __412806_412806;
   reg _412807_412807 ; 
   reg __412807_412807;
   reg _412808_412808 ; 
   reg __412808_412808;
   reg _412809_412809 ; 
   reg __412809_412809;
   reg _412810_412810 ; 
   reg __412810_412810;
   reg _412811_412811 ; 
   reg __412811_412811;
   reg _412812_412812 ; 
   reg __412812_412812;
   reg _412813_412813 ; 
   reg __412813_412813;
   reg _412814_412814 ; 
   reg __412814_412814;
   reg _412815_412815 ; 
   reg __412815_412815;
   reg _412816_412816 ; 
   reg __412816_412816;
   reg _412817_412817 ; 
   reg __412817_412817;
   reg _412818_412818 ; 
   reg __412818_412818;
   reg _412819_412819 ; 
   reg __412819_412819;
   reg _412820_412820 ; 
   reg __412820_412820;
   reg _412821_412821 ; 
   reg __412821_412821;
   reg _412822_412822 ; 
   reg __412822_412822;
   reg _412823_412823 ; 
   reg __412823_412823;
   reg _412824_412824 ; 
   reg __412824_412824;
   reg _412825_412825 ; 
   reg __412825_412825;
   reg _412826_412826 ; 
   reg __412826_412826;
   reg _412827_412827 ; 
   reg __412827_412827;
   reg _412828_412828 ; 
   reg __412828_412828;
   reg _412829_412829 ; 
   reg __412829_412829;
   reg _412830_412830 ; 
   reg __412830_412830;
   reg _412831_412831 ; 
   reg __412831_412831;
   reg _412832_412832 ; 
   reg __412832_412832;
   reg _412833_412833 ; 
   reg __412833_412833;
   reg _412834_412834 ; 
   reg __412834_412834;
   reg _412835_412835 ; 
   reg __412835_412835;
   reg _412836_412836 ; 
   reg __412836_412836;
   reg _412837_412837 ; 
   reg __412837_412837;
   reg _412838_412838 ; 
   reg __412838_412838;
   reg _412839_412839 ; 
   reg __412839_412839;
   reg _412840_412840 ; 
   reg __412840_412840;
   reg _412841_412841 ; 
   reg __412841_412841;
   reg _412842_412842 ; 
   reg __412842_412842;
   reg _412843_412843 ; 
   reg __412843_412843;
   reg _412844_412844 ; 
   reg __412844_412844;
   reg _412845_412845 ; 
   reg __412845_412845;
   reg _412846_412846 ; 
   reg __412846_412846;
   reg _412847_412847 ; 
   reg __412847_412847;
   reg _412848_412848 ; 
   reg __412848_412848;
   reg _412849_412849 ; 
   reg __412849_412849;
   reg _412850_412850 ; 
   reg __412850_412850;
   reg _412851_412851 ; 
   reg __412851_412851;
   reg _412852_412852 ; 
   reg __412852_412852;
   reg _412853_412853 ; 
   reg __412853_412853;
   reg _412854_412854 ; 
   reg __412854_412854;
   reg _412855_412855 ; 
   reg __412855_412855;
   reg _412856_412856 ; 
   reg __412856_412856;
   reg _412857_412857 ; 
   reg __412857_412857;
   reg _412858_412858 ; 
   reg __412858_412858;
   reg _412859_412859 ; 
   reg __412859_412859;
   reg _412860_412860 ; 
   reg __412860_412860;
   reg _412861_412861 ; 
   reg __412861_412861;
   reg _412862_412862 ; 
   reg __412862_412862;
   reg _412863_412863 ; 
   reg __412863_412863;
   reg _412864_412864 ; 
   reg __412864_412864;
   reg _412865_412865 ; 
   reg __412865_412865;
   reg _412866_412866 ; 
   reg __412866_412866;
   reg _412867_412867 ; 
   reg __412867_412867;
   reg _412868_412868 ; 
   reg __412868_412868;
   reg _412869_412869 ; 
   reg __412869_412869;
   reg _412870_412870 ; 
   reg __412870_412870;
   reg _412871_412871 ; 
   reg __412871_412871;
   reg _412872_412872 ; 
   reg __412872_412872;
   reg _412873_412873 ; 
   reg __412873_412873;
   reg _412874_412874 ; 
   reg __412874_412874;
   reg _412875_412875 ; 
   reg __412875_412875;
   reg _412876_412876 ; 
   reg __412876_412876;
   reg _412877_412877 ; 
   reg __412877_412877;
   reg _412878_412878 ; 
   reg __412878_412878;
   reg _412879_412879 ; 
   reg __412879_412879;
   reg _412880_412880 ; 
   reg __412880_412880;
   reg _412881_412881 ; 
   reg __412881_412881;
   reg _412882_412882 ; 
   reg __412882_412882;
   reg _412883_412883 ; 
   reg __412883_412883;
   reg _412884_412884 ; 
   reg __412884_412884;
   reg _412885_412885 ; 
   reg __412885_412885;
   reg _412886_412886 ; 
   reg __412886_412886;
   reg _412887_412887 ; 
   reg __412887_412887;
   reg _412888_412888 ; 
   reg __412888_412888;
   reg _412889_412889 ; 
   reg __412889_412889;
   reg _412890_412890 ; 
   reg __412890_412890;
   reg _412891_412891 ; 
   reg __412891_412891;
   reg _412892_412892 ; 
   reg __412892_412892;
   reg _412893_412893 ; 
   reg __412893_412893;
   reg _412894_412894 ; 
   reg __412894_412894;
   reg _412895_412895 ; 
   reg __412895_412895;
   reg _412896_412896 ; 
   reg __412896_412896;
   reg _412897_412897 ; 
   reg __412897_412897;
   reg _412898_412898 ; 
   reg __412898_412898;
   reg _412899_412899 ; 
   reg __412899_412899;
   reg _412900_412900 ; 
   reg __412900_412900;
   reg _412901_412901 ; 
   reg __412901_412901;
   reg _412902_412902 ; 
   reg __412902_412902;
   reg _412903_412903 ; 
   reg __412903_412903;
   reg _412904_412904 ; 
   reg __412904_412904;
   reg _412905_412905 ; 
   reg __412905_412905;
   reg _412906_412906 ; 
   reg __412906_412906;
   reg _412907_412907 ; 
   reg __412907_412907;
   reg _412908_412908 ; 
   reg __412908_412908;
   reg _412909_412909 ; 
   reg __412909_412909;
   reg _412910_412910 ; 
   reg __412910_412910;
   reg _412911_412911 ; 
   reg __412911_412911;
   reg _412912_412912 ; 
   reg __412912_412912;
   reg _412913_412913 ; 
   reg __412913_412913;
   reg _412914_412914 ; 
   reg __412914_412914;
   reg _412915_412915 ; 
   reg __412915_412915;
   reg _412916_412916 ; 
   reg __412916_412916;
   reg _412917_412917 ; 
   reg __412917_412917;
   reg _412918_412918 ; 
   reg __412918_412918;
   reg _412919_412919 ; 
   reg __412919_412919;
   reg _412920_412920 ; 
   reg __412920_412920;
   reg _412921_412921 ; 
   reg __412921_412921;
   reg _412922_412922 ; 
   reg __412922_412922;
   reg _412923_412923 ; 
   reg __412923_412923;
   reg _412924_412924 ; 
   reg __412924_412924;
   reg _412925_412925 ; 
   reg __412925_412925;
   reg _412926_412926 ; 
   reg __412926_412926;
   reg _412927_412927 ; 
   reg __412927_412927;
   reg _412928_412928 ; 
   reg __412928_412928;
   reg _412929_412929 ; 
   reg __412929_412929;
   reg _412930_412930 ; 
   reg __412930_412930;
   reg _412931_412931 ; 
   reg __412931_412931;
   reg _412932_412932 ; 
   reg __412932_412932;
   reg _412933_412933 ; 
   reg __412933_412933;
   reg _412934_412934 ; 
   reg __412934_412934;
   reg _412935_412935 ; 
   reg __412935_412935;
   reg _412936_412936 ; 
   reg __412936_412936;
   reg _412937_412937 ; 
   reg __412937_412937;
   reg _412938_412938 ; 
   reg __412938_412938;
   reg _412939_412939 ; 
   reg __412939_412939;
   reg _412940_412940 ; 
   reg __412940_412940;
   reg _412941_412941 ; 
   reg __412941_412941;
   reg _412942_412942 ; 
   reg __412942_412942;
   reg _412943_412943 ; 
   reg __412943_412943;
   reg _412944_412944 ; 
   reg __412944_412944;
   reg _412945_412945 ; 
   reg __412945_412945;
   reg _412946_412946 ; 
   reg __412946_412946;
   reg _412947_412947 ; 
   reg __412947_412947;
   reg _412948_412948 ; 
   reg __412948_412948;
   reg _412949_412949 ; 
   reg __412949_412949;
   reg _412950_412950 ; 
   reg __412950_412950;
   reg _412951_412951 ; 
   reg __412951_412951;
   reg _412952_412952 ; 
   reg __412952_412952;
   reg _412953_412953 ; 
   reg __412953_412953;
   reg _412954_412954 ; 
   reg __412954_412954;
   reg _412955_412955 ; 
   reg __412955_412955;
   reg _412956_412956 ; 
   reg __412956_412956;
   reg _412957_412957 ; 
   reg __412957_412957;
   reg _412958_412958 ; 
   reg __412958_412958;
   reg _412959_412959 ; 
   reg __412959_412959;
   reg _412960_412960 ; 
   reg __412960_412960;
   reg _412961_412961 ; 
   reg __412961_412961;
   reg _412962_412962 ; 
   reg __412962_412962;
   reg _412963_412963 ; 
   reg __412963_412963;
   reg _412964_412964 ; 
   reg __412964_412964;
   reg _412965_412965 ; 
   reg __412965_412965;
   reg _412966_412966 ; 
   reg __412966_412966;
   reg _412967_412967 ; 
   reg __412967_412967;
   reg _412968_412968 ; 
   reg __412968_412968;
   reg _412969_412969 ; 
   reg __412969_412969;
   reg _412970_412970 ; 
   reg __412970_412970;
   reg _412971_412971 ; 
   reg __412971_412971;
   reg _412972_412972 ; 
   reg __412972_412972;
   reg _412973_412973 ; 
   reg __412973_412973;
   reg _412974_412974 ; 
   reg __412974_412974;
   reg _412975_412975 ; 
   reg __412975_412975;
   reg _412976_412976 ; 
   reg __412976_412976;
   reg _412977_412977 ; 
   reg __412977_412977;
   reg _412978_412978 ; 
   reg __412978_412978;
   reg _412979_412979 ; 
   reg __412979_412979;
   reg _412980_412980 ; 
   reg __412980_412980;
   reg _412981_412981 ; 
   reg __412981_412981;
   reg _412982_412982 ; 
   reg __412982_412982;
   reg _412983_412983 ; 
   reg __412983_412983;
   reg _412984_412984 ; 
   reg __412984_412984;
   reg _412985_412985 ; 
   reg __412985_412985;
   reg _412986_412986 ; 
   reg __412986_412986;
   reg _412987_412987 ; 
   reg __412987_412987;
   reg _412988_412988 ; 
   reg __412988_412988;
   reg _412989_412989 ; 
   reg __412989_412989;
   reg _412990_412990 ; 
   reg __412990_412990;
   reg _412991_412991 ; 
   reg __412991_412991;
   reg _412992_412992 ; 
   reg __412992_412992;
   reg _412993_412993 ; 
   reg __412993_412993;
   reg _412994_412994 ; 
   reg __412994_412994;
   reg _412995_412995 ; 
   reg __412995_412995;
   reg _412996_412996 ; 
   reg __412996_412996;
   reg _412997_412997 ; 
   reg __412997_412997;
   reg _412998_412998 ; 
   reg __412998_412998;
   reg _412999_412999 ; 
   reg __412999_412999;
   reg _413000_413000 ; 
   reg __413000_413000;
   reg _413001_413001 ; 
   reg __413001_413001;
   reg _413002_413002 ; 
   reg __413002_413002;
   reg _413003_413003 ; 
   reg __413003_413003;
   reg _413004_413004 ; 
   reg __413004_413004;
   reg _413005_413005 ; 
   reg __413005_413005;
   reg _413006_413006 ; 
   reg __413006_413006;
   reg _413007_413007 ; 
   reg __413007_413007;
   reg _413008_413008 ; 
   reg __413008_413008;
   reg _413009_413009 ; 
   reg __413009_413009;
   reg _413010_413010 ; 
   reg __413010_413010;
   reg _413011_413011 ; 
   reg __413011_413011;
   reg _413012_413012 ; 
   reg __413012_413012;
   reg _413013_413013 ; 
   reg __413013_413013;
   reg _413014_413014 ; 
   reg __413014_413014;
   reg _413015_413015 ; 
   reg __413015_413015;
   reg _413016_413016 ; 
   reg __413016_413016;
   reg _413017_413017 ; 
   reg __413017_413017;
   reg _413018_413018 ; 
   reg __413018_413018;
   reg _413019_413019 ; 
   reg __413019_413019;
   reg _413020_413020 ; 
   reg __413020_413020;
   reg _413021_413021 ; 
   reg __413021_413021;
   reg _413022_413022 ; 
   reg __413022_413022;
   reg _413023_413023 ; 
   reg __413023_413023;
   reg _413024_413024 ; 
   reg __413024_413024;
   reg _413025_413025 ; 
   reg __413025_413025;
   reg _413026_413026 ; 
   reg __413026_413026;
   reg _413027_413027 ; 
   reg __413027_413027;
   reg _413028_413028 ; 
   reg __413028_413028;
   reg _413029_413029 ; 
   reg __413029_413029;
   reg _413030_413030 ; 
   reg __413030_413030;
   reg _413031_413031 ; 
   reg __413031_413031;
   reg _413032_413032 ; 
   reg __413032_413032;
   reg _413033_413033 ; 
   reg __413033_413033;
   reg _413034_413034 ; 
   reg __413034_413034;
   reg _413035_413035 ; 
   reg __413035_413035;
   reg _413036_413036 ; 
   reg __413036_413036;
   reg _413037_413037 ; 
   reg __413037_413037;
   reg _413038_413038 ; 
   reg __413038_413038;
   reg _413039_413039 ; 
   reg __413039_413039;
   reg _413040_413040 ; 
   reg __413040_413040;
   reg _413041_413041 ; 
   reg __413041_413041;
   reg _413042_413042 ; 
   reg __413042_413042;
   reg _413043_413043 ; 
   reg __413043_413043;
   reg _413044_413044 ; 
   reg __413044_413044;
   reg _413045_413045 ; 
   reg __413045_413045;
   reg _413046_413046 ; 
   reg __413046_413046;
   reg _413047_413047 ; 
   reg __413047_413047;
   reg _413048_413048 ; 
   reg __413048_413048;
   reg _413049_413049 ; 
   reg __413049_413049;
   reg _413050_413050 ; 
   reg __413050_413050;
   reg _413051_413051 ; 
   reg __413051_413051;
   reg _413052_413052 ; 
   reg __413052_413052;
   reg _413053_413053 ; 
   reg __413053_413053;
   reg _413054_413054 ; 
   reg __413054_413054;
   reg _413055_413055 ; 
   reg __413055_413055;
   reg _413056_413056 ; 
   reg __413056_413056;
   reg _413057_413057 ; 
   reg __413057_413057;
   reg _413058_413058 ; 
   reg __413058_413058;
   reg _413059_413059 ; 
   reg __413059_413059;
   reg _413060_413060 ; 
   reg __413060_413060;
   reg _413061_413061 ; 
   reg __413061_413061;
   reg _413062_413062 ; 
   reg __413062_413062;
   reg _413063_413063 ; 
   reg __413063_413063;
   reg _413064_413064 ; 
   reg __413064_413064;
   reg _413065_413065 ; 
   reg __413065_413065;
   reg _413066_413066 ; 
   reg __413066_413066;
   reg _413067_413067 ; 
   reg __413067_413067;
   reg _413068_413068 ; 
   reg __413068_413068;
   reg _413069_413069 ; 
   reg __413069_413069;
   reg _413070_413070 ; 
   reg __413070_413070;
   reg _413071_413071 ; 
   reg __413071_413071;
   reg _413072_413072 ; 
   reg __413072_413072;
   reg _413073_413073 ; 
   reg __413073_413073;
   reg _413074_413074 ; 
   reg __413074_413074;
   reg _413075_413075 ; 
   reg __413075_413075;
   reg _413076_413076 ; 
   reg __413076_413076;
   reg _413077_413077 ; 
   reg __413077_413077;
   reg _413078_413078 ; 
   reg __413078_413078;
   reg _413079_413079 ; 
   reg __413079_413079;
   reg _413080_413080 ; 
   reg __413080_413080;
   reg _413081_413081 ; 
   reg __413081_413081;
   reg _413082_413082 ; 
   reg __413082_413082;
   reg _413083_413083 ; 
   reg __413083_413083;
   reg _413084_413084 ; 
   reg __413084_413084;
   reg _413085_413085 ; 
   reg __413085_413085;
   reg _413086_413086 ; 
   reg __413086_413086;
   reg _413087_413087 ; 
   reg __413087_413087;
   reg _413088_413088 ; 
   reg __413088_413088;
   reg _413089_413089 ; 
   reg __413089_413089;
   reg _413090_413090 ; 
   reg __413090_413090;
   reg _413091_413091 ; 
   reg __413091_413091;
   reg _413092_413092 ; 
   reg __413092_413092;
   reg _413093_413093 ; 
   reg __413093_413093;
   reg _413094_413094 ; 
   reg __413094_413094;
   reg _413095_413095 ; 
   reg __413095_413095;
   reg _413096_413096 ; 
   reg __413096_413096;
   reg _413097_413097 ; 
   reg __413097_413097;
   reg _413098_413098 ; 
   reg __413098_413098;
   reg _413099_413099 ; 
   reg __413099_413099;
   reg _413100_413100 ; 
   reg __413100_413100;
   reg _413101_413101 ; 
   reg __413101_413101;
   reg _413102_413102 ; 
   reg __413102_413102;
   reg _413103_413103 ; 
   reg __413103_413103;
   reg _413104_413104 ; 
   reg __413104_413104;
   reg _413105_413105 ; 
   reg __413105_413105;
   reg _413106_413106 ; 
   reg __413106_413106;
   reg _413107_413107 ; 
   reg __413107_413107;
   reg _413108_413108 ; 
   reg __413108_413108;
   reg _413109_413109 ; 
   reg __413109_413109;
   reg _413110_413110 ; 
   reg __413110_413110;
   reg _413111_413111 ; 
   reg __413111_413111;
   reg _413112_413112 ; 
   reg __413112_413112;
   reg _413113_413113 ; 
   reg __413113_413113;
   reg _413114_413114 ; 
   reg __413114_413114;
   reg _413115_413115 ; 
   reg __413115_413115;
   reg _413116_413116 ; 
   reg __413116_413116;
   reg _413117_413117 ; 
   reg __413117_413117;
   reg _413118_413118 ; 
   reg __413118_413118;
   reg _413119_413119 ; 
   reg __413119_413119;
   reg _413120_413120 ; 
   reg __413120_413120;
   reg _413121_413121 ; 
   reg __413121_413121;
   reg _413122_413122 ; 
   reg __413122_413122;
   reg _413123_413123 ; 
   reg __413123_413123;
   reg _413124_413124 ; 
   reg __413124_413124;
   reg _413125_413125 ; 
   reg __413125_413125;
   reg _413126_413126 ; 
   reg __413126_413126;
   reg _413127_413127 ; 
   reg __413127_413127;
   reg _413128_413128 ; 
   reg __413128_413128;
   reg _413129_413129 ; 
   reg __413129_413129;
   reg _413130_413130 ; 
   reg __413130_413130;
   reg _413131_413131 ; 
   reg __413131_413131;
   reg _413132_413132 ; 
   reg __413132_413132;
   reg _413133_413133 ; 
   reg __413133_413133;
   reg _413134_413134 ; 
   reg __413134_413134;
   reg _413135_413135 ; 
   reg __413135_413135;
   reg _413136_413136 ; 
   reg __413136_413136;
   reg _413137_413137 ; 
   reg __413137_413137;
   reg _413138_413138 ; 
   reg __413138_413138;
   reg _413139_413139 ; 
   reg __413139_413139;
   reg _413140_413140 ; 
   reg __413140_413140;
   reg _413141_413141 ; 
   reg __413141_413141;
   reg _413142_413142 ; 
   reg __413142_413142;
   reg _413143_413143 ; 
   reg __413143_413143;
   reg _413144_413144 ; 
   reg __413144_413144;
   reg _413145_413145 ; 
   reg __413145_413145;
   reg _413146_413146 ; 
   reg __413146_413146;
   reg _413147_413147 ; 
   reg __413147_413147;
   reg _413148_413148 ; 
   reg __413148_413148;
   reg _413149_413149 ; 
   reg __413149_413149;
   reg _413150_413150 ; 
   reg __413150_413150;
   reg _413151_413151 ; 
   reg __413151_413151;
   reg _413152_413152 ; 
   reg __413152_413152;
   reg _413153_413153 ; 
   reg __413153_413153;
   reg _413154_413154 ; 
   reg __413154_413154;
   reg _413155_413155 ; 
   reg __413155_413155;
   reg _413156_413156 ; 
   reg __413156_413156;
   reg _413157_413157 ; 
   reg __413157_413157;
   reg _413158_413158 ; 
   reg __413158_413158;
   reg _413159_413159 ; 
   reg __413159_413159;
   reg _413160_413160 ; 
   reg __413160_413160;
   reg _413161_413161 ; 
   reg __413161_413161;
   reg _413162_413162 ; 
   reg __413162_413162;
   reg _413163_413163 ; 
   reg __413163_413163;
   reg _413164_413164 ; 
   reg __413164_413164;
   reg _413165_413165 ; 
   reg __413165_413165;
   reg _413166_413166 ; 
   reg __413166_413166;
   reg _413167_413167 ; 
   reg __413167_413167;
   reg _413168_413168 ; 
   reg __413168_413168;
   reg _413169_413169 ; 
   reg __413169_413169;
   reg _413170_413170 ; 
   reg __413170_413170;
   reg _413171_413171 ; 
   reg __413171_413171;
   reg _413172_413172 ; 
   reg __413172_413172;
   reg _413173_413173 ; 
   reg __413173_413173;
   reg _413174_413174 ; 
   reg __413174_413174;
   reg _413175_413175 ; 
   reg __413175_413175;
   reg _413176_413176 ; 
   reg __413176_413176;
   reg _413177_413177 ; 
   reg __413177_413177;
   reg _413178_413178 ; 
   reg __413178_413178;
   reg _413179_413179 ; 
   reg __413179_413179;
   reg _413180_413180 ; 
   reg __413180_413180;
   reg _413181_413181 ; 
   reg __413181_413181;
   reg _413182_413182 ; 
   reg __413182_413182;
   reg _413183_413183 ; 
   reg __413183_413183;
   reg _413184_413184 ; 
   reg __413184_413184;
   reg _413185_413185 ; 
   reg __413185_413185;
   reg _413186_413186 ; 
   reg __413186_413186;
   reg _413187_413187 ; 
   reg __413187_413187;
   reg _413188_413188 ; 
   reg __413188_413188;
   reg _413189_413189 ; 
   reg __413189_413189;
   reg _413190_413190 ; 
   reg __413190_413190;
   reg _413191_413191 ; 
   reg __413191_413191;
   reg _413192_413192 ; 
   reg __413192_413192;
   reg _413193_413193 ; 
   reg __413193_413193;
   reg _413194_413194 ; 
   reg __413194_413194;
   reg _413195_413195 ; 
   reg __413195_413195;
   reg _413196_413196 ; 
   reg __413196_413196;
   reg _413197_413197 ; 
   reg __413197_413197;
   reg _413198_413198 ; 
   reg __413198_413198;
   reg _413199_413199 ; 
   reg __413199_413199;
   reg _413200_413200 ; 
   reg __413200_413200;
   reg _413201_413201 ; 
   reg __413201_413201;
   reg _413202_413202 ; 
   reg __413202_413202;
   reg _413203_413203 ; 
   reg __413203_413203;
   reg _413204_413204 ; 
   reg __413204_413204;
   reg _413205_413205 ; 
   reg __413205_413205;
   reg _413206_413206 ; 
   reg __413206_413206;
   reg _413207_413207 ; 
   reg __413207_413207;
   reg _413208_413208 ; 
   reg __413208_413208;
   reg _413209_413209 ; 
   reg __413209_413209;
   reg _413210_413210 ; 
   reg __413210_413210;
   reg _413211_413211 ; 
   reg __413211_413211;
   reg _413212_413212 ; 
   reg __413212_413212;
   reg _413213_413213 ; 
   reg __413213_413213;
   reg _413214_413214 ; 
   reg __413214_413214;
   reg _413215_413215 ; 
   reg __413215_413215;
   reg _413216_413216 ; 
   reg __413216_413216;
   reg _413217_413217 ; 
   reg __413217_413217;
   reg _413218_413218 ; 
   reg __413218_413218;
   reg _413219_413219 ; 
   reg __413219_413219;
   reg _413220_413220 ; 
   reg __413220_413220;
   reg _413221_413221 ; 
   reg __413221_413221;
   reg _413222_413222 ; 
   reg __413222_413222;
   reg _413223_413223 ; 
   reg __413223_413223;
   reg _413224_413224 ; 
   reg __413224_413224;
   reg _413225_413225 ; 
   reg __413225_413225;
   reg _413226_413226 ; 
   reg __413226_413226;
   reg _413227_413227 ; 
   reg __413227_413227;
   reg _413228_413228 ; 
   reg __413228_413228;
   reg _413229_413229 ; 
   reg __413229_413229;
   reg _413230_413230 ; 
   reg __413230_413230;
   reg _413231_413231 ; 
   reg __413231_413231;
   reg _413232_413232 ; 
   reg __413232_413232;
   reg _413233_413233 ; 
   reg __413233_413233;
   reg _413234_413234 ; 
   reg __413234_413234;
   reg _413235_413235 ; 
   reg __413235_413235;
   reg _413236_413236 ; 
   reg __413236_413236;
   reg _413237_413237 ; 
   reg __413237_413237;
   reg _413238_413238 ; 
   reg __413238_413238;
   reg _413239_413239 ; 
   reg __413239_413239;
   reg _413240_413240 ; 
   reg __413240_413240;
   reg _413241_413241 ; 
   reg __413241_413241;
   reg _413242_413242 ; 
   reg __413242_413242;
   reg _413243_413243 ; 
   reg __413243_413243;
   reg _413244_413244 ; 
   reg __413244_413244;
   reg _413245_413245 ; 
   reg __413245_413245;
   reg _413246_413246 ; 
   reg __413246_413246;
   reg _413247_413247 ; 
   reg __413247_413247;
   reg _413248_413248 ; 
   reg __413248_413248;
   reg _413249_413249 ; 
   reg __413249_413249;
   reg _413250_413250 ; 
   reg __413250_413250;
   reg _413251_413251 ; 
   reg __413251_413251;
   reg _413252_413252 ; 
   reg __413252_413252;
   reg _413253_413253 ; 
   reg __413253_413253;
   reg _413254_413254 ; 
   reg __413254_413254;
   reg _413255_413255 ; 
   reg __413255_413255;
   reg _413256_413256 ; 
   reg __413256_413256;
   reg _413257_413257 ; 
   reg __413257_413257;
   reg _413258_413258 ; 
   reg __413258_413258;
   reg _413259_413259 ; 
   reg __413259_413259;
   reg _413260_413260 ; 
   reg __413260_413260;
   reg _413261_413261 ; 
   reg __413261_413261;
   reg _413262_413262 ; 
   reg __413262_413262;
   reg _413263_413263 ; 
   reg __413263_413263;
   reg _413264_413264 ; 
   reg __413264_413264;
   reg _413265_413265 ; 
   reg __413265_413265;
   reg _413266_413266 ; 
   reg __413266_413266;
   reg _413267_413267 ; 
   reg __413267_413267;
   reg _413268_413268 ; 
   reg __413268_413268;
   reg _413269_413269 ; 
   reg __413269_413269;
   reg _413270_413270 ; 
   reg __413270_413270;
   reg _413271_413271 ; 
   reg __413271_413271;
   reg _413272_413272 ; 
   reg __413272_413272;
   reg _413273_413273 ; 
   reg __413273_413273;
   reg _413274_413274 ; 
   reg __413274_413274;
   reg _413275_413275 ; 
   reg __413275_413275;
   reg _413276_413276 ; 
   reg __413276_413276;
   reg _413277_413277 ; 
   reg __413277_413277;
   reg _413278_413278 ; 
   reg __413278_413278;
   reg _413279_413279 ; 
   reg __413279_413279;
   reg _413280_413280 ; 
   reg __413280_413280;
   reg _413281_413281 ; 
   reg __413281_413281;
   reg _413282_413282 ; 
   reg __413282_413282;
   reg _413283_413283 ; 
   reg __413283_413283;
   reg _413284_413284 ; 
   reg __413284_413284;
   reg _413285_413285 ; 
   reg __413285_413285;
   reg _413286_413286 ; 
   reg __413286_413286;
   reg _413287_413287 ; 
   reg __413287_413287;
   reg _413288_413288 ; 
   reg __413288_413288;
   reg _413289_413289 ; 
   reg __413289_413289;
   reg _413290_413290 ; 
   reg __413290_413290;
   reg _413291_413291 ; 
   reg __413291_413291;
   reg _413292_413292 ; 
   reg __413292_413292;
   reg _413293_413293 ; 
   reg __413293_413293;
   reg _413294_413294 ; 
   reg __413294_413294;
   reg _413295_413295 ; 
   reg __413295_413295;
   reg _413296_413296 ; 
   reg __413296_413296;
   reg _413297_413297 ; 
   reg __413297_413297;
   reg _413298_413298 ; 
   reg __413298_413298;
   reg _413299_413299 ; 
   reg __413299_413299;
   reg _413300_413300 ; 
   reg __413300_413300;
   reg _413301_413301 ; 
   reg __413301_413301;
   reg _413302_413302 ; 
   reg __413302_413302;
   reg _413303_413303 ; 
   reg __413303_413303;
   reg _413304_413304 ; 
   reg __413304_413304;
   reg _413305_413305 ; 
   reg __413305_413305;
   reg _413306_413306 ; 
   reg __413306_413306;
   reg _413307_413307 ; 
   reg __413307_413307;
   reg _413308_413308 ; 
   reg __413308_413308;
   reg _413309_413309 ; 
   reg __413309_413309;
   reg _413310_413310 ; 
   reg __413310_413310;
   reg _413311_413311 ; 
   reg __413311_413311;
   reg _413312_413312 ; 
   reg __413312_413312;
   reg _413313_413313 ; 
   reg __413313_413313;
   reg _413314_413314 ; 
   reg __413314_413314;
   reg _413315_413315 ; 
   reg __413315_413315;
   reg _413316_413316 ; 
   reg __413316_413316;
   reg _413317_413317 ; 
   reg __413317_413317;
   reg _413318_413318 ; 
   reg __413318_413318;
   reg _413319_413319 ; 
   reg __413319_413319;
   reg _413320_413320 ; 
   reg __413320_413320;
   reg _413321_413321 ; 
   reg __413321_413321;
   reg _413322_413322 ; 
   reg __413322_413322;
   reg _413323_413323 ; 
   reg __413323_413323;
   reg _413324_413324 ; 
   reg __413324_413324;
   reg _413325_413325 ; 
   reg __413325_413325;
   reg _413326_413326 ; 
   reg __413326_413326;
   reg _413327_413327 ; 
   reg __413327_413327;
   reg _413328_413328 ; 
   reg __413328_413328;
   reg _413329_413329 ; 
   reg __413329_413329;
   reg _413330_413330 ; 
   reg __413330_413330;
   reg _413331_413331 ; 
   reg __413331_413331;
   reg _413332_413332 ; 
   reg __413332_413332;
   reg _413333_413333 ; 
   reg __413333_413333;
   reg _413334_413334 ; 
   reg __413334_413334;
   reg _413335_413335 ; 
   reg __413335_413335;
   reg _413336_413336 ; 
   reg __413336_413336;
   reg _413337_413337 ; 
   reg __413337_413337;
   reg _413338_413338 ; 
   reg __413338_413338;
   reg _413339_413339 ; 
   reg __413339_413339;
   reg _413340_413340 ; 
   reg __413340_413340;
   reg _413341_413341 ; 
   reg __413341_413341;
   reg _413342_413342 ; 
   reg __413342_413342;
   reg _413343_413343 ; 
   reg __413343_413343;
   reg _413344_413344 ; 
   reg __413344_413344;
   reg _413345_413345 ; 
   reg __413345_413345;
   reg _413346_413346 ; 
   reg __413346_413346;
   reg _413347_413347 ; 
   reg __413347_413347;
   reg _413348_413348 ; 
   reg __413348_413348;
   reg _413349_413349 ; 
   reg __413349_413349;
   reg _413350_413350 ; 
   reg __413350_413350;
   reg _413351_413351 ; 
   reg __413351_413351;
   reg _413352_413352 ; 
   reg __413352_413352;
   reg _413353_413353 ; 
   reg __413353_413353;
   reg _413354_413354 ; 
   reg __413354_413354;
   reg _413355_413355 ; 
   reg __413355_413355;
   reg _413356_413356 ; 
   reg __413356_413356;
   reg _413357_413357 ; 
   reg __413357_413357;
   reg _413358_413358 ; 
   reg __413358_413358;
   reg _413359_413359 ; 
   reg __413359_413359;
   reg _413360_413360 ; 
   reg __413360_413360;
   reg _413361_413361 ; 
   reg __413361_413361;
   reg _413362_413362 ; 
   reg __413362_413362;
   reg _413363_413363 ; 
   reg __413363_413363;
   reg _413364_413364 ; 
   reg __413364_413364;
   reg _413365_413365 ; 
   reg __413365_413365;
   reg _413366_413366 ; 
   reg __413366_413366;
   reg _413367_413367 ; 
   reg __413367_413367;
   reg _413368_413368 ; 
   reg __413368_413368;
   reg _413369_413369 ; 
   reg __413369_413369;
   reg _413370_413370 ; 
   reg __413370_413370;
   reg _413371_413371 ; 
   reg __413371_413371;
   reg _413372_413372 ; 
   reg __413372_413372;
   reg _413373_413373 ; 
   reg __413373_413373;
   reg _413374_413374 ; 
   reg __413374_413374;
   reg _413375_413375 ; 
   reg __413375_413375;
   reg _413376_413376 ; 
   reg __413376_413376;
   reg _413377_413377 ; 
   reg __413377_413377;
   reg _413378_413378 ; 
   reg __413378_413378;
   reg _413379_413379 ; 
   reg __413379_413379;
   reg _413380_413380 ; 
   reg __413380_413380;
   reg _413381_413381 ; 
   reg __413381_413381;
   reg _413382_413382 ; 
   reg __413382_413382;
   reg _413383_413383 ; 
   reg __413383_413383;
   reg _413384_413384 ; 
   reg __413384_413384;
   reg _413385_413385 ; 
   reg __413385_413385;
   reg _413386_413386 ; 
   reg __413386_413386;
   reg _413387_413387 ; 
   reg __413387_413387;
   reg _413388_413388 ; 
   reg __413388_413388;
   reg _413389_413389 ; 
   reg __413389_413389;
   reg _413390_413390 ; 
   reg __413390_413390;
   reg _413391_413391 ; 
   reg __413391_413391;
   reg _413392_413392 ; 
   reg __413392_413392;
   reg _413393_413393 ; 
   reg __413393_413393;
   reg _413394_413394 ; 
   reg __413394_413394;
   reg _413395_413395 ; 
   reg __413395_413395;
   reg _413396_413396 ; 
   reg __413396_413396;
   reg _413397_413397 ; 
   reg __413397_413397;
   reg _413398_413398 ; 
   reg __413398_413398;
   reg _413399_413399 ; 
   reg __413399_413399;
   reg _413400_413400 ; 
   reg __413400_413400;
   reg _413401_413401 ; 
   reg __413401_413401;
   reg _413402_413402 ; 
   reg __413402_413402;
   reg _413403_413403 ; 
   reg __413403_413403;
   reg _413404_413404 ; 
   reg __413404_413404;
   reg _413405_413405 ; 
   reg __413405_413405;
   reg _413406_413406 ; 
   reg __413406_413406;
   reg _413407_413407 ; 
   reg __413407_413407;
   reg _413408_413408 ; 
   reg __413408_413408;
   reg _413409_413409 ; 
   reg __413409_413409;
   reg _413410_413410 ; 
   reg __413410_413410;
   reg _413411_413411 ; 
   reg __413411_413411;
   reg _413412_413412 ; 
   reg __413412_413412;
   reg _413413_413413 ; 
   reg __413413_413413;
   reg _413414_413414 ; 
   reg __413414_413414;
   reg _413415_413415 ; 
   reg __413415_413415;
   reg _413416_413416 ; 
   reg __413416_413416;
   reg _413417_413417 ; 
   reg __413417_413417;
   reg _413418_413418 ; 
   reg __413418_413418;
   reg _413419_413419 ; 
   reg __413419_413419;
   reg _413420_413420 ; 
   reg __413420_413420;
   reg _413421_413421 ; 
   reg __413421_413421;
   reg _413422_413422 ; 
   reg __413422_413422;
   reg _413423_413423 ; 
   reg __413423_413423;
   reg _413424_413424 ; 
   reg __413424_413424;
   reg _413425_413425 ; 
   reg __413425_413425;
   reg _413426_413426 ; 
   reg __413426_413426;
   reg _413427_413427 ; 
   reg __413427_413427;
   reg _413428_413428 ; 
   reg __413428_413428;
   reg _413429_413429 ; 
   reg __413429_413429;
   reg _413430_413430 ; 
   reg __413430_413430;
   reg _413431_413431 ; 
   reg __413431_413431;
   reg _413432_413432 ; 
   reg __413432_413432;
   reg _413433_413433 ; 
   reg __413433_413433;
   reg _413434_413434 ; 
   reg __413434_413434;
   reg _413435_413435 ; 
   reg __413435_413435;
   reg _413436_413436 ; 
   reg __413436_413436;
   reg _413437_413437 ; 
   reg __413437_413437;
   reg _413438_413438 ; 
   reg __413438_413438;
   reg _413439_413439 ; 
   reg __413439_413439;
   reg _413440_413440 ; 
   reg __413440_413440;
   reg _413441_413441 ; 
   reg __413441_413441;
   reg _413442_413442 ; 
   reg __413442_413442;
   reg _413443_413443 ; 
   reg __413443_413443;
   reg _413444_413444 ; 
   reg __413444_413444;
   reg _413445_413445 ; 
   reg __413445_413445;
   reg _413446_413446 ; 
   reg __413446_413446;
   reg _413447_413447 ; 
   reg __413447_413447;
   reg _413448_413448 ; 
   reg __413448_413448;
   reg _413449_413449 ; 
   reg __413449_413449;
   reg _413450_413450 ; 
   reg __413450_413450;
   reg _413451_413451 ; 
   reg __413451_413451;
   reg _413452_413452 ; 
   reg __413452_413452;
   reg _413453_413453 ; 
   reg __413453_413453;
   reg _413454_413454 ; 
   reg __413454_413454;
   reg _413455_413455 ; 
   reg __413455_413455;
   reg _413456_413456 ; 
   reg __413456_413456;
   reg _413457_413457 ; 
   reg __413457_413457;
   reg _413458_413458 ; 
   reg __413458_413458;
   reg _413459_413459 ; 
   reg __413459_413459;
   reg _413460_413460 ; 
   reg __413460_413460;
   reg _413461_413461 ; 
   reg __413461_413461;
   reg _413462_413462 ; 
   reg __413462_413462;
   reg _413463_413463 ; 
   reg __413463_413463;
   reg _413464_413464 ; 
   reg __413464_413464;
   reg _413465_413465 ; 
   reg __413465_413465;
   reg _413466_413466 ; 
   reg __413466_413466;
   reg _413467_413467 ; 
   reg __413467_413467;
   reg _413468_413468 ; 
   reg __413468_413468;
   reg _413469_413469 ; 
   reg __413469_413469;
   reg _413470_413470 ; 
   reg __413470_413470;
   reg _413471_413471 ; 
   reg __413471_413471;
   reg _413472_413472 ; 
   reg __413472_413472;
   reg _413473_413473 ; 
   reg __413473_413473;
   reg _413474_413474 ; 
   reg __413474_413474;
   reg _413475_413475 ; 
   reg __413475_413475;
   reg _413476_413476 ; 
   reg __413476_413476;
   reg _413477_413477 ; 
   reg __413477_413477;
   reg _413478_413478 ; 
   reg __413478_413478;
   reg _413479_413479 ; 
   reg __413479_413479;
   reg _413480_413480 ; 
   reg __413480_413480;
   reg _413481_413481 ; 
   reg __413481_413481;
   reg _413482_413482 ; 
   reg __413482_413482;
   reg _413483_413483 ; 
   reg __413483_413483;
   reg _413484_413484 ; 
   reg __413484_413484;
   reg _413485_413485 ; 
   reg __413485_413485;
   reg _413486_413486 ; 
   reg __413486_413486;
   reg _413487_413487 ; 
   reg __413487_413487;
   reg _413488_413488 ; 
   reg __413488_413488;
   reg _413489_413489 ; 
   reg __413489_413489;
   reg _413490_413490 ; 
   reg __413490_413490;
   reg _413491_413491 ; 
   reg __413491_413491;
   reg _413492_413492 ; 
   reg __413492_413492;
   reg _413493_413493 ; 
   reg __413493_413493;
   reg _413494_413494 ; 
   reg __413494_413494;
   reg _413495_413495 ; 
   reg __413495_413495;
   reg _413496_413496 ; 
   reg __413496_413496;
   reg _413497_413497 ; 
   reg __413497_413497;
   reg _413498_413498 ; 
   reg __413498_413498;
   reg _413499_413499 ; 
   reg __413499_413499;
   reg _413500_413500 ; 
   reg __413500_413500;
   reg _413501_413501 ; 
   reg __413501_413501;
   reg _413502_413502 ; 
   reg __413502_413502;
   reg _413503_413503 ; 
   reg __413503_413503;
   reg _413504_413504 ; 
   reg __413504_413504;
   reg _413505_413505 ; 
   reg __413505_413505;
   reg _413506_413506 ; 
   reg __413506_413506;
   reg _413507_413507 ; 
   reg __413507_413507;
   reg _413508_413508 ; 
   reg __413508_413508;
   reg _413509_413509 ; 
   reg __413509_413509;
   reg _413510_413510 ; 
   reg __413510_413510;
   reg _413511_413511 ; 
   reg __413511_413511;
   reg _413512_413512 ; 
   reg __413512_413512;
   reg _413513_413513 ; 
   reg __413513_413513;
   reg _413514_413514 ; 
   reg __413514_413514;
   reg _413515_413515 ; 
   reg __413515_413515;
   reg _413516_413516 ; 
   reg __413516_413516;
   reg _413517_413517 ; 
   reg __413517_413517;
   reg _413518_413518 ; 
   reg __413518_413518;
   reg _413519_413519 ; 
   reg __413519_413519;
   reg _413520_413520 ; 
   reg __413520_413520;
   reg _413521_413521 ; 
   reg __413521_413521;
   reg _413522_413522 ; 
   reg __413522_413522;
   reg _413523_413523 ; 
   reg __413523_413523;
   reg _413524_413524 ; 
   reg __413524_413524;
   reg _413525_413525 ; 
   reg __413525_413525;
   reg _413526_413526 ; 
   reg __413526_413526;
   reg _413527_413527 ; 
   reg __413527_413527;
   reg _413528_413528 ; 
   reg __413528_413528;
   reg _413529_413529 ; 
   reg __413529_413529;
   reg _413530_413530 ; 
   reg __413530_413530;
   reg _413531_413531 ; 
   reg __413531_413531;
   reg _413532_413532 ; 
   reg __413532_413532;
   reg _413533_413533 ; 
   reg __413533_413533;
   reg _413534_413534 ; 
   reg __413534_413534;
   reg _413535_413535 ; 
   reg __413535_413535;
   reg _413536_413536 ; 
   reg __413536_413536;
   reg _413537_413537 ; 
   reg __413537_413537;
   reg _413538_413538 ; 
   reg __413538_413538;
   reg _413539_413539 ; 
   reg __413539_413539;
   reg _413540_413540 ; 
   reg __413540_413540;
   reg _413541_413541 ; 
   reg __413541_413541;
   reg _413542_413542 ; 
   reg __413542_413542;
   reg _413543_413543 ; 
   reg __413543_413543;
   reg _413544_413544 ; 
   reg __413544_413544;
   reg _413545_413545 ; 
   reg __413545_413545;
   reg _413546_413546 ; 
   reg __413546_413546;
   reg _413547_413547 ; 
   reg __413547_413547;
   reg _413548_413548 ; 
   reg __413548_413548;
   reg _413549_413549 ; 
   reg __413549_413549;
   reg _413550_413550 ; 
   reg __413550_413550;
   reg _413551_413551 ; 
   reg __413551_413551;
   reg _413552_413552 ; 
   reg __413552_413552;
   reg _413553_413553 ; 
   reg __413553_413553;
   reg _413554_413554 ; 
   reg __413554_413554;
   reg _413555_413555 ; 
   reg __413555_413555;
   reg _413556_413556 ; 
   reg __413556_413556;
   reg _413557_413557 ; 
   reg __413557_413557;
   reg _413558_413558 ; 
   reg __413558_413558;
   reg _413559_413559 ; 
   reg __413559_413559;
   reg _413560_413560 ; 
   reg __413560_413560;
   reg _413561_413561 ; 
   reg __413561_413561;
   reg _413562_413562 ; 
   reg __413562_413562;
   reg _413563_413563 ; 
   reg __413563_413563;
   reg _413564_413564 ; 
   reg __413564_413564;
   reg _413565_413565 ; 
   reg __413565_413565;
   reg _413566_413566 ; 
   reg __413566_413566;
   reg _413567_413567 ; 
   reg __413567_413567;
   reg _413568_413568 ; 
   reg __413568_413568;
   reg _413569_413569 ; 
   reg __413569_413569;
   reg _413570_413570 ; 
   reg __413570_413570;
   reg _413571_413571 ; 
   reg __413571_413571;
   reg _413572_413572 ; 
   reg __413572_413572;
   reg _413573_413573 ; 
   reg __413573_413573;
   reg _413574_413574 ; 
   reg __413574_413574;
   reg _413575_413575 ; 
   reg __413575_413575;
   reg _413576_413576 ; 
   reg __413576_413576;
   reg _413577_413577 ; 
   reg __413577_413577;
   reg _413578_413578 ; 
   reg __413578_413578;
   reg _413579_413579 ; 
   reg __413579_413579;
   reg _413580_413580 ; 
   reg __413580_413580;
   reg _413581_413581 ; 
   reg __413581_413581;
   reg _413582_413582 ; 
   reg __413582_413582;
   reg _413583_413583 ; 
   reg __413583_413583;
   reg _413584_413584 ; 
   reg __413584_413584;
   reg _413585_413585 ; 
   reg __413585_413585;
   reg _413586_413586 ; 
   reg __413586_413586;
   reg _413587_413587 ; 
   reg __413587_413587;
   reg _413588_413588 ; 
   reg __413588_413588;
   reg _413589_413589 ; 
   reg __413589_413589;
   reg _413590_413590 ; 
   reg __413590_413590;
   reg _413591_413591 ; 
   reg __413591_413591;
   reg _413592_413592 ; 
   reg __413592_413592;
   reg _413593_413593 ; 
   reg __413593_413593;
   reg _413594_413594 ; 
   reg __413594_413594;
   reg _413595_413595 ; 
   reg __413595_413595;
   reg _413596_413596 ; 
   reg __413596_413596;
   reg _413597_413597 ; 
   reg __413597_413597;
   reg _413598_413598 ; 
   reg __413598_413598;
   reg _413599_413599 ; 
   reg __413599_413599;
   reg _413600_413600 ; 
   reg __413600_413600;
   reg _413601_413601 ; 
   reg __413601_413601;
   reg _413602_413602 ; 
   reg __413602_413602;
   reg _413603_413603 ; 
   reg __413603_413603;
   reg _413604_413604 ; 
   reg __413604_413604;
   reg _413605_413605 ; 
   reg __413605_413605;
   reg _413606_413606 ; 
   reg __413606_413606;
   reg _413607_413607 ; 
   reg __413607_413607;
   reg _413608_413608 ; 
   reg __413608_413608;
   reg _413609_413609 ; 
   reg __413609_413609;
   reg _413610_413610 ; 
   reg __413610_413610;
   reg _413611_413611 ; 
   reg __413611_413611;
   reg _413612_413612 ; 
   reg __413612_413612;
   reg _413613_413613 ; 
   reg __413613_413613;
   reg _413614_413614 ; 
   reg __413614_413614;
   reg _413615_413615 ; 
   reg __413615_413615;
   reg _413616_413616 ; 
   reg __413616_413616;
   reg _413617_413617 ; 
   reg __413617_413617;
   reg _413618_413618 ; 
   reg __413618_413618;
   reg _413619_413619 ; 
   reg __413619_413619;
   reg _413620_413620 ; 
   reg __413620_413620;
   reg _413621_413621 ; 
   reg __413621_413621;
   reg _413622_413622 ; 
   reg __413622_413622;
   reg _413623_413623 ; 
   reg __413623_413623;
   reg _413624_413624 ; 
   reg __413624_413624;
   reg _413625_413625 ; 
   reg __413625_413625;
   reg _413626_413626 ; 
   reg __413626_413626;
   reg _413627_413627 ; 
   reg __413627_413627;
   reg _413628_413628 ; 
   reg __413628_413628;
   reg _413629_413629 ; 
   reg __413629_413629;
   reg _413630_413630 ; 
   reg __413630_413630;
   reg _413631_413631 ; 
   reg __413631_413631;
   reg _413632_413632 ; 
   reg __413632_413632;
   reg _413633_413633 ; 
   reg __413633_413633;
   reg _413634_413634 ; 
   reg __413634_413634;
   reg _413635_413635 ; 
   reg __413635_413635;
   reg _413636_413636 ; 
   reg __413636_413636;
   reg _413637_413637 ; 
   reg __413637_413637;
   reg _413638_413638 ; 
   reg __413638_413638;
   reg _413639_413639 ; 
   reg __413639_413639;
   reg _413640_413640 ; 
   reg __413640_413640;
   reg _413641_413641 ; 
   reg __413641_413641;
   reg _413642_413642 ; 
   reg __413642_413642;
   reg _413643_413643 ; 
   reg __413643_413643;
   reg _413644_413644 ; 
   reg __413644_413644;
   reg _413645_413645 ; 
   reg __413645_413645;
   reg _413646_413646 ; 
   reg __413646_413646;
   reg _413647_413647 ; 
   reg __413647_413647;
   reg _413648_413648 ; 
   reg __413648_413648;
   reg _413649_413649 ; 
   reg __413649_413649;
   reg _413650_413650 ; 
   reg __413650_413650;
   reg _413651_413651 ; 
   reg __413651_413651;
   reg _413652_413652 ; 
   reg __413652_413652;
   reg _413653_413653 ; 
   reg __413653_413653;
   reg _413654_413654 ; 
   reg __413654_413654;
   reg _413655_413655 ; 
   reg __413655_413655;
   reg _413656_413656 ; 
   reg __413656_413656;
   reg _413657_413657 ; 
   reg __413657_413657;
   reg _413658_413658 ; 
   reg __413658_413658;
   reg _413659_413659 ; 
   reg __413659_413659;
   reg _413660_413660 ; 
   reg __413660_413660;
   reg _413661_413661 ; 
   reg __413661_413661;
   reg _413662_413662 ; 
   reg __413662_413662;
   reg _413663_413663 ; 
   reg __413663_413663;
   reg _413664_413664 ; 
   reg __413664_413664;
   reg _413665_413665 ; 
   reg __413665_413665;
   reg _413666_413666 ; 
   reg __413666_413666;
   reg _413667_413667 ; 
   reg __413667_413667;
   reg _413668_413668 ; 
   reg __413668_413668;
   reg _413669_413669 ; 
   reg __413669_413669;
   reg _413670_413670 ; 
   reg __413670_413670;
   reg _413671_413671 ; 
   reg __413671_413671;
   reg _413672_413672 ; 
   reg __413672_413672;
   reg _413673_413673 ; 
   reg __413673_413673;
   reg _413674_413674 ; 
   reg __413674_413674;
   reg _413675_413675 ; 
   reg __413675_413675;
   reg _413676_413676 ; 
   reg __413676_413676;
   reg _413677_413677 ; 
   reg __413677_413677;
   reg _413678_413678 ; 
   reg __413678_413678;
   reg _413679_413679 ; 
   reg __413679_413679;
   reg _413680_413680 ; 
   reg __413680_413680;
   reg _413681_413681 ; 
   reg __413681_413681;
   reg _413682_413682 ; 
   reg __413682_413682;
   reg _413683_413683 ; 
   reg __413683_413683;
   reg _413684_413684 ; 
   reg __413684_413684;
   reg _413685_413685 ; 
   reg __413685_413685;
   reg _413686_413686 ; 
   reg __413686_413686;
   reg _413687_413687 ; 
   reg __413687_413687;
   reg _413688_413688 ; 
   reg __413688_413688;
   reg _413689_413689 ; 
   reg __413689_413689;
   reg _413690_413690 ; 
   reg __413690_413690;
   reg _413691_413691 ; 
   reg __413691_413691;
   reg _413692_413692 ; 
   reg __413692_413692;
   reg _413693_413693 ; 
   reg __413693_413693;
   reg _413694_413694 ; 
   reg __413694_413694;
   reg _413695_413695 ; 
   reg __413695_413695;
   reg _413696_413696 ; 
   reg __413696_413696;
   reg _413697_413697 ; 
   reg __413697_413697;
   reg _413698_413698 ; 
   reg __413698_413698;
   reg _413699_413699 ; 
   reg __413699_413699;
   reg _413700_413700 ; 
   reg __413700_413700;
   reg _413701_413701 ; 
   reg __413701_413701;
   reg _413702_413702 ; 
   reg __413702_413702;
   reg _413703_413703 ; 
   reg __413703_413703;
   reg _413704_413704 ; 
   reg __413704_413704;
   reg _413705_413705 ; 
   reg __413705_413705;
   reg _413706_413706 ; 
   reg __413706_413706;
   reg _413707_413707 ; 
   reg __413707_413707;
   reg _413708_413708 ; 
   reg __413708_413708;
   reg _413709_413709 ; 
   reg __413709_413709;
   reg _413710_413710 ; 
   reg __413710_413710;
   reg _413711_413711 ; 
   reg __413711_413711;
   reg _413712_413712 ; 
   reg __413712_413712;
   reg _413713_413713 ; 
   reg __413713_413713;
   reg _413714_413714 ; 
   reg __413714_413714;
   reg _413715_413715 ; 
   reg __413715_413715;
   reg _413716_413716 ; 
   reg __413716_413716;
   reg _413717_413717 ; 
   reg __413717_413717;
   reg _413718_413718 ; 
   reg __413718_413718;
   reg _413719_413719 ; 
   reg __413719_413719;
   reg _413720_413720 ; 
   reg __413720_413720;
   reg _413721_413721 ; 
   reg __413721_413721;
   reg _413722_413722 ; 
   reg __413722_413722;
   reg _413723_413723 ; 
   reg __413723_413723;
   reg _413724_413724 ; 
   reg __413724_413724;
   reg _413725_413725 ; 
   reg __413725_413725;
   reg _413726_413726 ; 
   reg __413726_413726;
   reg _413727_413727 ; 
   reg __413727_413727;
   reg _413728_413728 ; 
   reg __413728_413728;
   reg _413729_413729 ; 
   reg __413729_413729;
   reg _413730_413730 ; 
   reg __413730_413730;
   reg _413731_413731 ; 
   reg __413731_413731;
   reg _413732_413732 ; 
   reg __413732_413732;
   reg _413733_413733 ; 
   reg __413733_413733;
   reg _413734_413734 ; 
   reg __413734_413734;
   reg _413735_413735 ; 
   reg __413735_413735;
   reg _413736_413736 ; 
   reg __413736_413736;
   reg _413737_413737 ; 
   reg __413737_413737;
   reg _413738_413738 ; 
   reg __413738_413738;
   reg _413739_413739 ; 
   reg __413739_413739;
   reg _413740_413740 ; 
   reg __413740_413740;
   reg _413741_413741 ; 
   reg __413741_413741;
   reg _413742_413742 ; 
   reg __413742_413742;
   reg _413743_413743 ; 
   reg __413743_413743;
   reg _413744_413744 ; 
   reg __413744_413744;
   reg _413745_413745 ; 
   reg __413745_413745;
   reg _413746_413746 ; 
   reg __413746_413746;
   reg _413747_413747 ; 
   reg __413747_413747;
   reg _413748_413748 ; 
   reg __413748_413748;
   reg _413749_413749 ; 
   reg __413749_413749;
   reg _413750_413750 ; 
   reg __413750_413750;
   reg _413751_413751 ; 
   reg __413751_413751;
   reg _413752_413752 ; 
   reg __413752_413752;
   reg _413753_413753 ; 
   reg __413753_413753;
   reg _413754_413754 ; 
   reg __413754_413754;
   reg _413755_413755 ; 
   reg __413755_413755;
   reg _413756_413756 ; 
   reg __413756_413756;
   reg _413757_413757 ; 
   reg __413757_413757;
   reg _413758_413758 ; 
   reg __413758_413758;
   reg _413759_413759 ; 
   reg __413759_413759;
   reg _413760_413760 ; 
   reg __413760_413760;
   reg _413761_413761 ; 
   reg __413761_413761;
   reg _413762_413762 ; 
   reg __413762_413762;
   reg _413763_413763 ; 
   reg __413763_413763;
   reg _413764_413764 ; 
   reg __413764_413764;
   reg _413765_413765 ; 
   reg __413765_413765;
   reg _413766_413766 ; 
   reg __413766_413766;
   reg _413767_413767 ; 
   reg __413767_413767;
   reg _413768_413768 ; 
   reg __413768_413768;
   reg _413769_413769 ; 
   reg __413769_413769;
   reg _413770_413770 ; 
   reg __413770_413770;
   reg _413771_413771 ; 
   reg __413771_413771;
   reg _413772_413772 ; 
   reg __413772_413772;
   reg _413773_413773 ; 
   reg __413773_413773;
   reg _413774_413774 ; 
   reg __413774_413774;
   reg _413775_413775 ; 
   reg __413775_413775;
   reg _413776_413776 ; 
   reg __413776_413776;
   reg _413777_413777 ; 
   reg __413777_413777;
   reg _413778_413778 ; 
   reg __413778_413778;
   reg _413779_413779 ; 
   reg __413779_413779;
   reg _413780_413780 ; 
   reg __413780_413780;
   reg _413781_413781 ; 
   reg __413781_413781;
   reg _413782_413782 ; 
   reg __413782_413782;
   reg _413783_413783 ; 
   reg __413783_413783;
   reg _413784_413784 ; 
   reg __413784_413784;
   reg _413785_413785 ; 
   reg __413785_413785;
   reg _413786_413786 ; 
   reg __413786_413786;
   reg _413787_413787 ; 
   reg __413787_413787;
   reg _413788_413788 ; 
   reg __413788_413788;
   reg _413789_413789 ; 
   reg __413789_413789;
   reg _413790_413790 ; 
   reg __413790_413790;
   reg _413791_413791 ; 
   reg __413791_413791;
   reg _413792_413792 ; 
   reg __413792_413792;
   reg _413793_413793 ; 
   reg __413793_413793;
   reg _413794_413794 ; 
   reg __413794_413794;
   reg _413795_413795 ; 
   reg __413795_413795;
   reg _413796_413796 ; 
   reg __413796_413796;
   reg _413797_413797 ; 
   reg __413797_413797;
   reg _413798_413798 ; 
   reg __413798_413798;
   reg _413799_413799 ; 
   reg __413799_413799;
   reg _413800_413800 ; 
   reg __413800_413800;
   reg _413801_413801 ; 
   reg __413801_413801;
   reg _413802_413802 ; 
   reg __413802_413802;
   reg _413803_413803 ; 
   reg __413803_413803;
   reg _413804_413804 ; 
   reg __413804_413804;
   reg _413805_413805 ; 
   reg __413805_413805;
   reg _413806_413806 ; 
   reg __413806_413806;
   reg _413807_413807 ; 
   reg __413807_413807;
   reg _413808_413808 ; 
   reg __413808_413808;
   reg _413809_413809 ; 
   reg __413809_413809;
   reg _413810_413810 ; 
   reg __413810_413810;
   reg _413811_413811 ; 
   reg __413811_413811;
   reg _413812_413812 ; 
   reg __413812_413812;
   reg _413813_413813 ; 
   reg __413813_413813;
   reg _413814_413814 ; 
   reg __413814_413814;
   reg _413815_413815 ; 
   reg __413815_413815;
   reg _413816_413816 ; 
   reg __413816_413816;
   reg _413817_413817 ; 
   reg __413817_413817;
   reg _413818_413818 ; 
   reg __413818_413818;
   reg _413819_413819 ; 
   reg __413819_413819;
   reg _413820_413820 ; 
   reg __413820_413820;
   reg _413821_413821 ; 
   reg __413821_413821;
   reg _413822_413822 ; 
   reg __413822_413822;
   reg _413823_413823 ; 
   reg __413823_413823;
   reg _413824_413824 ; 
   reg __413824_413824;
   reg _413825_413825 ; 
   reg __413825_413825;
   reg _413826_413826 ; 
   reg __413826_413826;
   reg _413827_413827 ; 
   reg __413827_413827;
   reg _413828_413828 ; 
   reg __413828_413828;
   reg _413829_413829 ; 
   reg __413829_413829;
   reg _413830_413830 ; 
   reg __413830_413830;
   reg _413831_413831 ; 
   reg __413831_413831;
   reg _413832_413832 ; 
   reg __413832_413832;
   reg _413833_413833 ; 
   reg __413833_413833;
   reg _413834_413834 ; 
   reg __413834_413834;
   reg _413835_413835 ; 
   reg __413835_413835;
   reg _413836_413836 ; 
   reg __413836_413836;
   reg _413837_413837 ; 
   reg __413837_413837;
   reg _413838_413838 ; 
   reg __413838_413838;
   reg _413839_413839 ; 
   reg __413839_413839;
   reg _413840_413840 ; 
   reg __413840_413840;
   reg _413841_413841 ; 
   reg __413841_413841;
   reg _413842_413842 ; 
   reg __413842_413842;
   reg _413843_413843 ; 
   reg __413843_413843;
   reg _413844_413844 ; 
   reg __413844_413844;
   reg _413845_413845 ; 
   reg __413845_413845;
   reg _413846_413846 ; 
   reg __413846_413846;
   reg _413847_413847 ; 
   reg __413847_413847;
   reg _413848_413848 ; 
   reg __413848_413848;
   reg _413849_413849 ; 
   reg __413849_413849;
   reg _413850_413850 ; 
   reg __413850_413850;
   reg _413851_413851 ; 
   reg __413851_413851;
   reg _413852_413852 ; 
   reg __413852_413852;
   reg _413853_413853 ; 
   reg __413853_413853;
   reg _413854_413854 ; 
   reg __413854_413854;
   reg _413855_413855 ; 
   reg __413855_413855;
   reg _413856_413856 ; 
   reg __413856_413856;
   reg _413857_413857 ; 
   reg __413857_413857;
   reg _413858_413858 ; 
   reg __413858_413858;
   reg _413859_413859 ; 
   reg __413859_413859;
   reg _413860_413860 ; 
   reg __413860_413860;
   reg _413861_413861 ; 
   reg __413861_413861;
   reg _413862_413862 ; 
   reg __413862_413862;
   reg _413863_413863 ; 
   reg __413863_413863;
   reg _413864_413864 ; 
   reg __413864_413864;
   reg _413865_413865 ; 
   reg __413865_413865;
   reg _413866_413866 ; 
   reg __413866_413866;
   reg _413867_413867 ; 
   reg __413867_413867;
   reg _413868_413868 ; 
   reg __413868_413868;
   reg _413869_413869 ; 
   reg __413869_413869;
   reg _413870_413870 ; 
   reg __413870_413870;
   reg _413871_413871 ; 
   reg __413871_413871;
   reg _413872_413872 ; 
   reg __413872_413872;
   reg _413873_413873 ; 
   reg __413873_413873;
   reg _413874_413874 ; 
   reg __413874_413874;
   reg _413875_413875 ; 
   reg __413875_413875;
   reg _413876_413876 ; 
   reg __413876_413876;
   reg _413877_413877 ; 
   reg __413877_413877;
   reg _413878_413878 ; 
   reg __413878_413878;
   reg _413879_413879 ; 
   reg __413879_413879;
   reg _413880_413880 ; 
   reg __413880_413880;
   reg _413881_413881 ; 
   reg __413881_413881;
   reg _413882_413882 ; 
   reg __413882_413882;
   reg _413883_413883 ; 
   reg __413883_413883;
   reg _413884_413884 ; 
   reg __413884_413884;
   reg _413885_413885 ; 
   reg __413885_413885;
   reg _413886_413886 ; 
   reg __413886_413886;
   reg _413887_413887 ; 
   reg __413887_413887;
   reg _413888_413888 ; 
   reg __413888_413888;
   reg _413889_413889 ; 
   reg __413889_413889;
   reg _413890_413890 ; 
   reg __413890_413890;
   reg _413891_413891 ; 
   reg __413891_413891;
   reg _413892_413892 ; 
   reg __413892_413892;
   reg _413893_413893 ; 
   reg __413893_413893;
   reg _413894_413894 ; 
   reg __413894_413894;
   reg _413895_413895 ; 
   reg __413895_413895;
   reg _413896_413896 ; 
   reg __413896_413896;
   reg _413897_413897 ; 
   reg __413897_413897;
   reg _413898_413898 ; 
   reg __413898_413898;
   reg _413899_413899 ; 
   reg __413899_413899;
   reg _413900_413900 ; 
   reg __413900_413900;
   reg _413901_413901 ; 
   reg __413901_413901;
   reg _413902_413902 ; 
   reg __413902_413902;
   reg _413903_413903 ; 
   reg __413903_413903;
   reg _413904_413904 ; 
   reg __413904_413904;
   reg _413905_413905 ; 
   reg __413905_413905;
   reg _413906_413906 ; 
   reg __413906_413906;
   reg _413907_413907 ; 
   reg __413907_413907;
   reg _413908_413908 ; 
   reg __413908_413908;
   reg _413909_413909 ; 
   reg __413909_413909;
   reg _413910_413910 ; 
   reg __413910_413910;
   reg _413911_413911 ; 
   reg __413911_413911;
   reg _413912_413912 ; 
   reg __413912_413912;
   reg _413913_413913 ; 
   reg __413913_413913;
   reg _413914_413914 ; 
   reg __413914_413914;
   reg _413915_413915 ; 
   reg __413915_413915;
   reg _413916_413916 ; 
   reg __413916_413916;
   reg _413917_413917 ; 
   reg __413917_413917;
   reg _413918_413918 ; 
   reg __413918_413918;
   reg _413919_413919 ; 
   reg __413919_413919;
   reg _413920_413920 ; 
   reg __413920_413920;
   reg _413921_413921 ; 
   reg __413921_413921;
   reg _413922_413922 ; 
   reg __413922_413922;
   reg _413923_413923 ; 
   reg __413923_413923;
   reg _413924_413924 ; 
   reg __413924_413924;
   reg _413925_413925 ; 
   reg __413925_413925;
   reg _413926_413926 ; 
   reg __413926_413926;
   reg _413927_413927 ; 
   reg __413927_413927;
   reg _413928_413928 ; 
   reg __413928_413928;
   reg _413929_413929 ; 
   reg __413929_413929;
   reg _413930_413930 ; 
   reg __413930_413930;
   reg _413931_413931 ; 
   reg __413931_413931;
   reg _413932_413932 ; 
   reg __413932_413932;
   reg _413933_413933 ; 
   reg __413933_413933;
   reg _413934_413934 ; 
   reg __413934_413934;
   reg _413935_413935 ; 
   reg __413935_413935;
   reg _413936_413936 ; 
   reg __413936_413936;
   reg _413937_413937 ; 
   reg __413937_413937;
   reg _413938_413938 ; 
   reg __413938_413938;
   reg _413939_413939 ; 
   reg __413939_413939;
   reg _413940_413940 ; 
   reg __413940_413940;
   reg _413941_413941 ; 
   reg __413941_413941;
   reg _413942_413942 ; 
   reg __413942_413942;
   reg _413943_413943 ; 
   reg __413943_413943;
   reg _413944_413944 ; 
   reg __413944_413944;
   reg _413945_413945 ; 
   reg __413945_413945;
   reg _413946_413946 ; 
   reg __413946_413946;
   reg _413947_413947 ; 
   reg __413947_413947;
   reg _413948_413948 ; 
   reg __413948_413948;
   reg _413949_413949 ; 
   reg __413949_413949;
   reg _413950_413950 ; 
   reg __413950_413950;
   reg _413951_413951 ; 
   reg __413951_413951;
   reg _413952_413952 ; 
   reg __413952_413952;
   reg _413953_413953 ; 
   reg __413953_413953;
   reg _413954_413954 ; 
   reg __413954_413954;
   reg _413955_413955 ; 
   reg __413955_413955;
   reg _413956_413956 ; 
   reg __413956_413956;
   reg _413957_413957 ; 
   reg __413957_413957;
   reg _413958_413958 ; 
   reg __413958_413958;
   reg _413959_413959 ; 
   reg __413959_413959;
   reg _413960_413960 ; 
   reg __413960_413960;
   reg _413961_413961 ; 
   reg __413961_413961;
   reg _413962_413962 ; 
   reg __413962_413962;
   reg _413963_413963 ; 
   reg __413963_413963;
   reg _413964_413964 ; 
   reg __413964_413964;
   reg _413965_413965 ; 
   reg __413965_413965;
   reg _413966_413966 ; 
   reg __413966_413966;
   reg _413967_413967 ; 
   reg __413967_413967;
   reg _413968_413968 ; 
   reg __413968_413968;
   reg _413969_413969 ; 
   reg __413969_413969;
   reg _413970_413970 ; 
   reg __413970_413970;
   reg _413971_413971 ; 
   reg __413971_413971;
   reg _413972_413972 ; 
   reg __413972_413972;
   reg _413973_413973 ; 
   reg __413973_413973;
   reg _413974_413974 ; 
   reg __413974_413974;
   reg _413975_413975 ; 
   reg __413975_413975;
   reg _413976_413976 ; 
   reg __413976_413976;
   reg _413977_413977 ; 
   reg __413977_413977;
   reg _413978_413978 ; 
   reg __413978_413978;
   reg _413979_413979 ; 
   reg __413979_413979;
   reg _413980_413980 ; 
   reg __413980_413980;
   reg _413981_413981 ; 
   reg __413981_413981;
   reg _413982_413982 ; 
   reg __413982_413982;
   reg _413983_413983 ; 
   reg __413983_413983;
   reg _413984_413984 ; 
   reg __413984_413984;
   reg _413985_413985 ; 
   reg __413985_413985;
   reg _413986_413986 ; 
   reg __413986_413986;
   reg _413987_413987 ; 
   reg __413987_413987;
   reg _413988_413988 ; 
   reg __413988_413988;
   reg _413989_413989 ; 
   reg __413989_413989;
   reg _413990_413990 ; 
   reg __413990_413990;
   reg _413991_413991 ; 
   reg __413991_413991;
   reg _413992_413992 ; 
   reg __413992_413992;
   reg _413993_413993 ; 
   reg __413993_413993;
   reg _413994_413994 ; 
   reg __413994_413994;
   reg _413995_413995 ; 
   reg __413995_413995;
   reg _413996_413996 ; 
   reg __413996_413996;
   reg _413997_413997 ; 
   reg __413997_413997;
   reg _413998_413998 ; 
   reg __413998_413998;
   reg _413999_413999 ; 
   reg __413999_413999;
   reg _414000_414000 ; 
   reg __414000_414000;
   reg _414001_414001 ; 
   reg __414001_414001;
   reg _414002_414002 ; 
   reg __414002_414002;
   reg _414003_414003 ; 
   reg __414003_414003;
   reg _414004_414004 ; 
   reg __414004_414004;
   reg _414005_414005 ; 
   reg __414005_414005;
   reg _414006_414006 ; 
   reg __414006_414006;
   reg _414007_414007 ; 
   reg __414007_414007;
   reg _414008_414008 ; 
   reg __414008_414008;
   reg _414009_414009 ; 
   reg __414009_414009;
   reg _414010_414010 ; 
   reg __414010_414010;
   reg _414011_414011 ; 
   reg __414011_414011;
   reg _414012_414012 ; 
   reg __414012_414012;
   reg _414013_414013 ; 
   reg __414013_414013;
   reg _414014_414014 ; 
   reg __414014_414014;
   reg _414015_414015 ; 
   reg __414015_414015;
   reg _414016_414016 ; 
   reg __414016_414016;
   reg _414017_414017 ; 
   reg __414017_414017;
   reg _414018_414018 ; 
   reg __414018_414018;
   reg _414019_414019 ; 
   reg __414019_414019;
   reg _414020_414020 ; 
   reg __414020_414020;
   reg _414021_414021 ; 
   reg __414021_414021;
   reg _414022_414022 ; 
   reg __414022_414022;
   reg _414023_414023 ; 
   reg __414023_414023;
   reg _414024_414024 ; 
   reg __414024_414024;
   reg _414025_414025 ; 
   reg __414025_414025;
   reg _414026_414026 ; 
   reg __414026_414026;
   reg _414027_414027 ; 
   reg __414027_414027;
   reg _414028_414028 ; 
   reg __414028_414028;
   reg _414029_414029 ; 
   reg __414029_414029;
   reg _414030_414030 ; 
   reg __414030_414030;
   reg _414031_414031 ; 
   reg __414031_414031;
   reg _414032_414032 ; 
   reg __414032_414032;
   reg _414033_414033 ; 
   reg __414033_414033;
   reg _414034_414034 ; 
   reg __414034_414034;
   reg _414035_414035 ; 
   reg __414035_414035;
   reg _414036_414036 ; 
   reg __414036_414036;
   reg _414037_414037 ; 
   reg __414037_414037;
   reg _414038_414038 ; 
   reg __414038_414038;
   reg _414039_414039 ; 
   reg __414039_414039;
   reg _414040_414040 ; 
   reg __414040_414040;
   reg _414041_414041 ; 
   reg __414041_414041;
   reg _414042_414042 ; 
   reg __414042_414042;
   reg _414043_414043 ; 
   reg __414043_414043;
   reg _414044_414044 ; 
   reg __414044_414044;
   reg _414045_414045 ; 
   reg __414045_414045;
   reg _414046_414046 ; 
   reg __414046_414046;
   reg _414047_414047 ; 
   reg __414047_414047;
   reg _414048_414048 ; 
   reg __414048_414048;
   reg _414049_414049 ; 
   reg __414049_414049;
   reg _414050_414050 ; 
   reg __414050_414050;
   reg _414051_414051 ; 
   reg __414051_414051;
   reg _414052_414052 ; 
   reg __414052_414052;
   reg _414053_414053 ; 
   reg __414053_414053;
   reg _414054_414054 ; 
   reg __414054_414054;
   reg _414055_414055 ; 
   reg __414055_414055;
   reg _414056_414056 ; 
   reg __414056_414056;
   reg _414057_414057 ; 
   reg __414057_414057;
   reg _414058_414058 ; 
   reg __414058_414058;
   reg _414059_414059 ; 
   reg __414059_414059;
   reg _414060_414060 ; 
   reg __414060_414060;
   reg _414061_414061 ; 
   reg __414061_414061;
   reg _414062_414062 ; 
   reg __414062_414062;
   reg _414063_414063 ; 
   reg __414063_414063;
   reg _414064_414064 ; 
   reg __414064_414064;
   reg _414065_414065 ; 
   reg __414065_414065;
   reg _414066_414066 ; 
   reg __414066_414066;
   reg _414067_414067 ; 
   reg __414067_414067;
   reg _414068_414068 ; 
   reg __414068_414068;
   reg _414069_414069 ; 
   reg __414069_414069;
   reg _414070_414070 ; 
   reg __414070_414070;
   reg _414071_414071 ; 
   reg __414071_414071;
   reg _414072_414072 ; 
   reg __414072_414072;
   reg _414073_414073 ; 
   reg __414073_414073;
   reg _414074_414074 ; 
   reg __414074_414074;
   reg _414075_414075 ; 
   reg __414075_414075;
   reg _414076_414076 ; 
   reg __414076_414076;
   reg _414077_414077 ; 
   reg __414077_414077;
   reg _414078_414078 ; 
   reg __414078_414078;
   reg _414079_414079 ; 
   reg __414079_414079;
   reg _414080_414080 ; 
   reg __414080_414080;
   reg _414081_414081 ; 
   reg __414081_414081;
   reg _414082_414082 ; 
   reg __414082_414082;
   reg _414083_414083 ; 
   reg __414083_414083;
   reg _414084_414084 ; 
   reg __414084_414084;
   reg _414085_414085 ; 
   reg __414085_414085;
   reg _414086_414086 ; 
   reg __414086_414086;
   reg _414087_414087 ; 
   reg __414087_414087;
   reg _414088_414088 ; 
   reg __414088_414088;
   reg _414089_414089 ; 
   reg __414089_414089;
   reg _414090_414090 ; 
   reg __414090_414090;
   reg _414091_414091 ; 
   reg __414091_414091;
   reg _414092_414092 ; 
   reg __414092_414092;
   reg _414093_414093 ; 
   reg __414093_414093;
   reg _414094_414094 ; 
   reg __414094_414094;
   reg _414095_414095 ; 
   reg __414095_414095;
   reg _414096_414096 ; 
   reg __414096_414096;
   reg _414097_414097 ; 
   reg __414097_414097;
   reg _414098_414098 ; 
   reg __414098_414098;
   reg _414099_414099 ; 
   reg __414099_414099;
   reg _414100_414100 ; 
   reg __414100_414100;
   reg _414101_414101 ; 
   reg __414101_414101;
   reg _414102_414102 ; 
   reg __414102_414102;
   reg _414103_414103 ; 
   reg __414103_414103;
   reg _414104_414104 ; 
   reg __414104_414104;
   reg _414105_414105 ; 
   reg __414105_414105;
   reg _414106_414106 ; 
   reg __414106_414106;
   reg _414107_414107 ; 
   reg __414107_414107;
   reg _414108_414108 ; 
   reg __414108_414108;
   reg _414109_414109 ; 
   reg __414109_414109;
   reg _414110_414110 ; 
   reg __414110_414110;
   reg _414111_414111 ; 
   reg __414111_414111;
   reg _414112_414112 ; 
   reg __414112_414112;
   reg _414113_414113 ; 
   reg __414113_414113;
   reg _414114_414114 ; 
   reg __414114_414114;
   reg _414115_414115 ; 
   reg __414115_414115;
   reg _414116_414116 ; 
   reg __414116_414116;
   reg _414117_414117 ; 
   reg __414117_414117;
   reg _414118_414118 ; 
   reg __414118_414118;
   reg _414119_414119 ; 
   reg __414119_414119;
   reg _414120_414120 ; 
   reg __414120_414120;
   reg _414121_414121 ; 
   reg __414121_414121;
   reg _414122_414122 ; 
   reg __414122_414122;
   reg _414123_414123 ; 
   reg __414123_414123;
   reg _414124_414124 ; 
   reg __414124_414124;
   reg _414125_414125 ; 
   reg __414125_414125;
   reg _414126_414126 ; 
   reg __414126_414126;
   reg _414127_414127 ; 
   reg __414127_414127;
   reg _414128_414128 ; 
   reg __414128_414128;
   reg _414129_414129 ; 
   reg __414129_414129;
   reg _414130_414130 ; 
   reg __414130_414130;
   reg _414131_414131 ; 
   reg __414131_414131;
   reg _414132_414132 ; 
   reg __414132_414132;
   reg _414133_414133 ; 
   reg __414133_414133;
   reg _414134_414134 ; 
   reg __414134_414134;
   reg _414135_414135 ; 
   reg __414135_414135;
   reg _414136_414136 ; 
   reg __414136_414136;
   reg _414137_414137 ; 
   reg __414137_414137;
   reg _414138_414138 ; 
   reg __414138_414138;
   reg _414139_414139 ; 
   reg __414139_414139;
   reg _414140_414140 ; 
   reg __414140_414140;
   reg _414141_414141 ; 
   reg __414141_414141;
   reg _414142_414142 ; 
   reg __414142_414142;
   reg _414143_414143 ; 
   reg __414143_414143;
   reg _414144_414144 ; 
   reg __414144_414144;
   reg _414145_414145 ; 
   reg __414145_414145;
   reg _414146_414146 ; 
   reg __414146_414146;
   reg _414147_414147 ; 
   reg __414147_414147;
   reg _414148_414148 ; 
   reg __414148_414148;
   reg _414149_414149 ; 
   reg __414149_414149;
   reg _414150_414150 ; 
   reg __414150_414150;
   reg _414151_414151 ; 
   reg __414151_414151;
   reg _414152_414152 ; 
   reg __414152_414152;
   reg _414153_414153 ; 
   reg __414153_414153;
   reg _414154_414154 ; 
   reg __414154_414154;
   reg _414155_414155 ; 
   reg __414155_414155;
   reg _414156_414156 ; 
   reg __414156_414156;
   reg _414157_414157 ; 
   reg __414157_414157;
   reg _414158_414158 ; 
   reg __414158_414158;
   reg _414159_414159 ; 
   reg __414159_414159;
   reg _414160_414160 ; 
   reg __414160_414160;
   reg _414161_414161 ; 
   reg __414161_414161;
   reg _414162_414162 ; 
   reg __414162_414162;
   reg _414163_414163 ; 
   reg __414163_414163;
   reg _414164_414164 ; 
   reg __414164_414164;
   reg _414165_414165 ; 
   reg __414165_414165;
   reg _414166_414166 ; 
   reg __414166_414166;
   reg _414167_414167 ; 
   reg __414167_414167;
   reg _414168_414168 ; 
   reg __414168_414168;
   reg _414169_414169 ; 
   reg __414169_414169;
   reg _414170_414170 ; 
   reg __414170_414170;
   reg _414171_414171 ; 
   reg __414171_414171;
   reg _414172_414172 ; 
   reg __414172_414172;
   reg _414173_414173 ; 
   reg __414173_414173;
   reg _414174_414174 ; 
   reg __414174_414174;
   reg _414175_414175 ; 
   reg __414175_414175;
   reg _414176_414176 ; 
   reg __414176_414176;
   reg _414177_414177 ; 
   reg __414177_414177;
   reg _414178_414178 ; 
   reg __414178_414178;
   reg _414179_414179 ; 
   reg __414179_414179;
   reg _414180_414180 ; 
   reg __414180_414180;
   reg _414181_414181 ; 
   reg __414181_414181;
   reg _414182_414182 ; 
   reg __414182_414182;
   reg _414183_414183 ; 
   reg __414183_414183;
   reg _414184_414184 ; 
   reg __414184_414184;
   reg _414185_414185 ; 
   reg __414185_414185;
   reg _414186_414186 ; 
   reg __414186_414186;
   reg _414187_414187 ; 
   reg __414187_414187;
   reg _414188_414188 ; 
   reg __414188_414188;
   reg _414189_414189 ; 
   reg __414189_414189;
   reg _414190_414190 ; 
   reg __414190_414190;
   reg _414191_414191 ; 
   reg __414191_414191;
   reg _414192_414192 ; 
   reg __414192_414192;
   reg _414193_414193 ; 
   reg __414193_414193;
   reg _414194_414194 ; 
   reg __414194_414194;
   reg _414195_414195 ; 
   reg __414195_414195;
   reg _414196_414196 ; 
   reg __414196_414196;
   reg _414197_414197 ; 
   reg __414197_414197;
   reg _414198_414198 ; 
   reg __414198_414198;
   reg _414199_414199 ; 
   reg __414199_414199;
   reg _414200_414200 ; 
   reg __414200_414200;
   reg _414201_414201 ; 
   reg __414201_414201;
   reg _414202_414202 ; 
   reg __414202_414202;
   reg _414203_414203 ; 
   reg __414203_414203;
   reg _414204_414204 ; 
   reg __414204_414204;
   reg _414205_414205 ; 
   reg __414205_414205;
   reg _414206_414206 ; 
   reg __414206_414206;
   reg _414207_414207 ; 
   reg __414207_414207;
   reg _414208_414208 ; 
   reg __414208_414208;
   reg _414209_414209 ; 
   reg __414209_414209;
   reg _414210_414210 ; 
   reg __414210_414210;
   reg _414211_414211 ; 
   reg __414211_414211;
   reg _414212_414212 ; 
   reg __414212_414212;
   reg _414213_414213 ; 
   reg __414213_414213;
   reg _414214_414214 ; 
   reg __414214_414214;
   reg _414215_414215 ; 
   reg __414215_414215;
   reg _414216_414216 ; 
   reg __414216_414216;
   reg _414217_414217 ; 
   reg __414217_414217;
   reg _414218_414218 ; 
   reg __414218_414218;
   reg _414219_414219 ; 
   reg __414219_414219;
   reg _414220_414220 ; 
   reg __414220_414220;
   reg _414221_414221 ; 
   reg __414221_414221;
   reg _414222_414222 ; 
   reg __414222_414222;
   reg _414223_414223 ; 
   reg __414223_414223;
   reg _414224_414224 ; 
   reg __414224_414224;
   reg _414225_414225 ; 
   reg __414225_414225;
   reg _414226_414226 ; 
   reg __414226_414226;
   reg _414227_414227 ; 
   reg __414227_414227;
   reg _414228_414228 ; 
   reg __414228_414228;
   reg _414229_414229 ; 
   reg __414229_414229;
   reg _414230_414230 ; 
   reg __414230_414230;
   reg _414231_414231 ; 
   reg __414231_414231;
   reg _414232_414232 ; 
   reg __414232_414232;
   reg _414233_414233 ; 
   reg __414233_414233;
   reg _414234_414234 ; 
   reg __414234_414234;
   reg _414235_414235 ; 
   reg __414235_414235;
   reg _414236_414236 ; 
   reg __414236_414236;
   reg _414237_414237 ; 
   reg __414237_414237;
   reg _414238_414238 ; 
   reg __414238_414238;
   reg _414239_414239 ; 
   reg __414239_414239;
   reg _414240_414240 ; 
   reg __414240_414240;
   reg _414241_414241 ; 
   reg __414241_414241;
   reg _414242_414242 ; 
   reg __414242_414242;
   reg _414243_414243 ; 
   reg __414243_414243;
   reg _414244_414244 ; 
   reg __414244_414244;
   reg _414245_414245 ; 
   reg __414245_414245;
   reg _414246_414246 ; 
   reg __414246_414246;
   reg _414247_414247 ; 
   reg __414247_414247;
   reg _414248_414248 ; 
   reg __414248_414248;
   reg _414249_414249 ; 
   reg __414249_414249;
   reg _414250_414250 ; 
   reg __414250_414250;
   reg _414251_414251 ; 
   reg __414251_414251;
   reg _414252_414252 ; 
   reg __414252_414252;
   reg _414253_414253 ; 
   reg __414253_414253;
   reg _414254_414254 ; 
   reg __414254_414254;
   reg _414255_414255 ; 
   reg __414255_414255;
   reg _414256_414256 ; 
   reg __414256_414256;
   reg _414257_414257 ; 
   reg __414257_414257;
   reg _414258_414258 ; 
   reg __414258_414258;
   reg _414259_414259 ; 
   reg __414259_414259;
   reg _414260_414260 ; 
   reg __414260_414260;
   reg _414261_414261 ; 
   reg __414261_414261;
   reg _414262_414262 ; 
   reg __414262_414262;
   reg _414263_414263 ; 
   reg __414263_414263;
   reg _414264_414264 ; 
   reg __414264_414264;
   reg _414265_414265 ; 
   reg __414265_414265;
   reg _414266_414266 ; 
   reg __414266_414266;
   reg _414267_414267 ; 
   reg __414267_414267;
   reg _414268_414268 ; 
   reg __414268_414268;
   reg _414269_414269 ; 
   reg __414269_414269;
   reg _414270_414270 ; 
   reg __414270_414270;
   reg _414271_414271 ; 
   reg __414271_414271;
   reg _414272_414272 ; 
   reg __414272_414272;
   reg _414273_414273 ; 
   reg __414273_414273;
   reg _414274_414274 ; 
   reg __414274_414274;
   reg _414275_414275 ; 
   reg __414275_414275;
   reg _414276_414276 ; 
   reg __414276_414276;
   reg _414277_414277 ; 
   reg __414277_414277;
   reg _414278_414278 ; 
   reg __414278_414278;
   reg _414279_414279 ; 
   reg __414279_414279;
   reg _414280_414280 ; 
   reg __414280_414280;
   reg _414281_414281 ; 
   reg __414281_414281;
   reg _414282_414282 ; 
   reg __414282_414282;
   reg _414283_414283 ; 
   reg __414283_414283;
   reg _414284_414284 ; 
   reg __414284_414284;
   reg _414285_414285 ; 
   reg __414285_414285;
   reg _414286_414286 ; 
   reg __414286_414286;
   reg _414287_414287 ; 
   reg __414287_414287;
   reg _414288_414288 ; 
   reg __414288_414288;
   reg _414289_414289 ; 
   reg __414289_414289;
   reg _414290_414290 ; 
   reg __414290_414290;
   reg _414291_414291 ; 
   reg __414291_414291;
   reg _414292_414292 ; 
   reg __414292_414292;
   reg _414293_414293 ; 
   reg __414293_414293;
   reg _414294_414294 ; 
   reg __414294_414294;
   reg _414295_414295 ; 
   reg __414295_414295;
   reg _414296_414296 ; 
   reg __414296_414296;
   reg _414297_414297 ; 
   reg __414297_414297;
   reg _414298_414298 ; 
   reg __414298_414298;
   reg _414299_414299 ; 
   reg __414299_414299;
   reg _414300_414300 ; 
   reg __414300_414300;
   reg _414301_414301 ; 
   reg __414301_414301;
   reg _414302_414302 ; 
   reg __414302_414302;
   reg _414303_414303 ; 
   reg __414303_414303;
   reg _414304_414304 ; 
   reg __414304_414304;
   reg _414305_414305 ; 
   reg __414305_414305;
   reg _414306_414306 ; 
   reg __414306_414306;
   reg _414307_414307 ; 
   reg __414307_414307;
   reg _414308_414308 ; 
   reg __414308_414308;
   reg _414309_414309 ; 
   reg __414309_414309;
   reg _414310_414310 ; 
   reg __414310_414310;
   reg _414311_414311 ; 
   reg __414311_414311;
   reg _414312_414312 ; 
   reg __414312_414312;
   reg _414313_414313 ; 
   reg __414313_414313;
   reg _414314_414314 ; 
   reg __414314_414314;
   reg _414315_414315 ; 
   reg __414315_414315;
   reg _414316_414316 ; 
   reg __414316_414316;
   reg _414317_414317 ; 
   reg __414317_414317;
   reg _414318_414318 ; 
   reg __414318_414318;
   reg _414319_414319 ; 
   reg __414319_414319;
   reg _414320_414320 ; 
   reg __414320_414320;
   reg _414321_414321 ; 
   reg __414321_414321;
   reg _414322_414322 ; 
   reg __414322_414322;
   reg _414323_414323 ; 
   reg __414323_414323;
   reg _414324_414324 ; 
   reg __414324_414324;
   reg _414325_414325 ; 
   reg __414325_414325;
   reg _414326_414326 ; 
   reg __414326_414326;
   reg _414327_414327 ; 
   reg __414327_414327;
   reg _414328_414328 ; 
   reg __414328_414328;
   reg _414329_414329 ; 
   reg __414329_414329;
   reg _414330_414330 ; 
   reg __414330_414330;
   reg _414331_414331 ; 
   reg __414331_414331;
   reg _414332_414332 ; 
   reg __414332_414332;
   reg _414333_414333 ; 
   reg __414333_414333;
   reg _414334_414334 ; 
   reg __414334_414334;
   reg _414335_414335 ; 
   reg __414335_414335;
   reg _414336_414336 ; 
   reg __414336_414336;
   reg _414337_414337 ; 
   reg __414337_414337;
   reg _414338_414338 ; 
   reg __414338_414338;
   reg _414339_414339 ; 
   reg __414339_414339;
   reg _414340_414340 ; 
   reg __414340_414340;
   reg _414341_414341 ; 
   reg __414341_414341;
   reg _414342_414342 ; 
   reg __414342_414342;
   reg _414343_414343 ; 
   reg __414343_414343;
   reg _414344_414344 ; 
   reg __414344_414344;
   reg _414345_414345 ; 
   reg __414345_414345;
   reg _414346_414346 ; 
   reg __414346_414346;
   reg _414347_414347 ; 
   reg __414347_414347;
   reg _414348_414348 ; 
   reg __414348_414348;
   reg _414349_414349 ; 
   reg __414349_414349;
   reg _414350_414350 ; 
   reg __414350_414350;
   reg _414351_414351 ; 
   reg __414351_414351;
   reg _414352_414352 ; 
   reg __414352_414352;
   reg _414353_414353 ; 
   reg __414353_414353;
   reg _414354_414354 ; 
   reg __414354_414354;
   reg _414355_414355 ; 
   reg __414355_414355;
   reg _414356_414356 ; 
   reg __414356_414356;
   reg _414357_414357 ; 
   reg __414357_414357;
   reg _414358_414358 ; 
   reg __414358_414358;
   reg _414359_414359 ; 
   reg __414359_414359;
   reg _414360_414360 ; 
   reg __414360_414360;
   reg _414361_414361 ; 
   reg __414361_414361;
   reg _414362_414362 ; 
   reg __414362_414362;
   reg _414363_414363 ; 
   reg __414363_414363;
   reg _414364_414364 ; 
   reg __414364_414364;
   reg _414365_414365 ; 
   reg __414365_414365;
   reg _414366_414366 ; 
   reg __414366_414366;
   reg _414367_414367 ; 
   reg __414367_414367;
   reg _414368_414368 ; 
   reg __414368_414368;
   reg _414369_414369 ; 
   reg __414369_414369;
   reg _414370_414370 ; 
   reg __414370_414370;
   reg _414371_414371 ; 
   reg __414371_414371;
   reg _414372_414372 ; 
   reg __414372_414372;
   reg _414373_414373 ; 
   reg __414373_414373;
   reg _414374_414374 ; 
   reg __414374_414374;
   reg _414375_414375 ; 
   reg __414375_414375;
   reg _414376_414376 ; 
   reg __414376_414376;
   reg _414377_414377 ; 
   reg __414377_414377;
   reg _414378_414378 ; 
   reg __414378_414378;
   reg _414379_414379 ; 
   reg __414379_414379;
   reg _414380_414380 ; 
   reg __414380_414380;
   reg _414381_414381 ; 
   reg __414381_414381;
   reg _414382_414382 ; 
   reg __414382_414382;
   reg _414383_414383 ; 
   reg __414383_414383;
   reg _414384_414384 ; 
   reg __414384_414384;
   reg _414385_414385 ; 
   reg __414385_414385;
   reg _414386_414386 ; 
   reg __414386_414386;
   reg _414387_414387 ; 
   reg __414387_414387;
   reg _414388_414388 ; 
   reg __414388_414388;
   reg _414389_414389 ; 
   reg __414389_414389;
   reg _414390_414390 ; 
   reg __414390_414390;
   reg _414391_414391 ; 
   reg __414391_414391;
   reg _414392_414392 ; 
   reg __414392_414392;
   reg _414393_414393 ; 
   reg __414393_414393;
   reg _414394_414394 ; 
   reg __414394_414394;
   reg _414395_414395 ; 
   reg __414395_414395;
   reg _414396_414396 ; 
   reg __414396_414396;
   reg _414397_414397 ; 
   reg __414397_414397;
   reg _414398_414398 ; 
   reg __414398_414398;
   reg _414399_414399 ; 
   reg __414399_414399;
   reg _414400_414400 ; 
   reg __414400_414400;
   reg _414401_414401 ; 
   reg __414401_414401;
   reg _414402_414402 ; 
   reg __414402_414402;
   reg _414403_414403 ; 
   reg __414403_414403;
   reg _414404_414404 ; 
   reg __414404_414404;
   reg _414405_414405 ; 
   reg __414405_414405;
   reg _414406_414406 ; 
   reg __414406_414406;
   reg _414407_414407 ; 
   reg __414407_414407;
   reg _414408_414408 ; 
   reg __414408_414408;
   reg _414409_414409 ; 
   reg __414409_414409;
   reg _414410_414410 ; 
   reg __414410_414410;
   reg _414411_414411 ; 
   reg __414411_414411;
   reg _414412_414412 ; 
   reg __414412_414412;
   reg _414413_414413 ; 
   reg __414413_414413;
   reg _414414_414414 ; 
   reg __414414_414414;
   reg _414415_414415 ; 
   reg __414415_414415;
   reg _414416_414416 ; 
   reg __414416_414416;
   reg _414417_414417 ; 
   reg __414417_414417;
   reg _414418_414418 ; 
   reg __414418_414418;
   reg _414419_414419 ; 
   reg __414419_414419;
   reg _414420_414420 ; 
   reg __414420_414420;
   reg _414421_414421 ; 
   reg __414421_414421;
   reg _414422_414422 ; 
   reg __414422_414422;
   reg _414423_414423 ; 
   reg __414423_414423;
   reg _414424_414424 ; 
   reg __414424_414424;
   reg _414425_414425 ; 
   reg __414425_414425;
   reg _414426_414426 ; 
   reg __414426_414426;
   reg _414427_414427 ; 
   reg __414427_414427;
   reg _414428_414428 ; 
   reg __414428_414428;
   reg _414429_414429 ; 
   reg __414429_414429;
   reg _414430_414430 ; 
   reg __414430_414430;
   reg _414431_414431 ; 
   reg __414431_414431;
   reg _414432_414432 ; 
   reg __414432_414432;
   reg _414433_414433 ; 
   reg __414433_414433;
   reg _414434_414434 ; 
   reg __414434_414434;
   reg _414435_414435 ; 
   reg __414435_414435;
   reg _414436_414436 ; 
   reg __414436_414436;
   reg _414437_414437 ; 
   reg __414437_414437;
   reg _414438_414438 ; 
   reg __414438_414438;
   reg _414439_414439 ; 
   reg __414439_414439;
   reg _414440_414440 ; 
   reg __414440_414440;
   reg _414441_414441 ; 
   reg __414441_414441;
   reg _414442_414442 ; 
   reg __414442_414442;
   reg _414443_414443 ; 
   reg __414443_414443;
   reg _414444_414444 ; 
   reg __414444_414444;
   reg _414445_414445 ; 
   reg __414445_414445;
   reg _414446_414446 ; 
   reg __414446_414446;
   reg _414447_414447 ; 
   reg __414447_414447;
   reg _414448_414448 ; 
   reg __414448_414448;
   reg _414449_414449 ; 
   reg __414449_414449;
   reg _414450_414450 ; 
   reg __414450_414450;
   reg _414451_414451 ; 
   reg __414451_414451;
   reg _414452_414452 ; 
   reg __414452_414452;
   reg _414453_414453 ; 
   reg __414453_414453;
   reg _414454_414454 ; 
   reg __414454_414454;
   reg _414455_414455 ; 
   reg __414455_414455;
   reg _414456_414456 ; 
   reg __414456_414456;
   reg _414457_414457 ; 
   reg __414457_414457;
   reg _414458_414458 ; 
   reg __414458_414458;
   reg _414459_414459 ; 
   reg __414459_414459;
   reg _414460_414460 ; 
   reg __414460_414460;
   reg _414461_414461 ; 
   reg __414461_414461;
   reg _414462_414462 ; 
   reg __414462_414462;
   reg _414463_414463 ; 
   reg __414463_414463;
   reg _414464_414464 ; 
   reg __414464_414464;
   reg _414465_414465 ; 
   reg __414465_414465;
   reg _414466_414466 ; 
   reg __414466_414466;
   reg _414467_414467 ; 
   reg __414467_414467;
   reg _414468_414468 ; 
   reg __414468_414468;
   reg _414469_414469 ; 
   reg __414469_414469;
   reg _414470_414470 ; 
   reg __414470_414470;
   reg _414471_414471 ; 
   reg __414471_414471;
   reg _414472_414472 ; 
   reg __414472_414472;
   reg _414473_414473 ; 
   reg __414473_414473;
   reg _414474_414474 ; 
   reg __414474_414474;
   reg _414475_414475 ; 
   reg __414475_414475;
   reg _414476_414476 ; 
   reg __414476_414476;
   reg _414477_414477 ; 
   reg __414477_414477;
   reg _414478_414478 ; 
   reg __414478_414478;
   reg _414479_414479 ; 
   reg __414479_414479;
   reg _414480_414480 ; 
   reg __414480_414480;
   reg _414481_414481 ; 
   reg __414481_414481;
   reg _414482_414482 ; 
   reg __414482_414482;
   reg _414483_414483 ; 
   reg __414483_414483;
   reg _414484_414484 ; 
   reg __414484_414484;
   reg _414485_414485 ; 
   reg __414485_414485;
   reg _414486_414486 ; 
   reg __414486_414486;
   reg _414487_414487 ; 
   reg __414487_414487;
   reg _414488_414488 ; 
   reg __414488_414488;
   reg _414489_414489 ; 
   reg __414489_414489;
   reg _414490_414490 ; 
   reg __414490_414490;
   reg _414491_414491 ; 
   reg __414491_414491;
   reg _414492_414492 ; 
   reg __414492_414492;
   reg _414493_414493 ; 
   reg __414493_414493;
   reg _414494_414494 ; 
   reg __414494_414494;
endmodule
