`include "defines.v"

module g1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 219
  output [1 - 1:0] ar_sa0_s10;
  f1 f10(.ar_sa0_s10(ar_sa0_s10));
  `include "g1.logic.vh"
endmodule

