// Test type: Binary Numbers - with spaces
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=5 'b01101;
endmodule
