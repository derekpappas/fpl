//test type : module_or_generate_item ::= parameter_override
//vparser rule name : 
//author : Codrin
module test_0260;
 (* in1 = 1, out2 *)
 defparam a.delay = 3;
endmodule
