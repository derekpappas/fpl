//test type : module_or_generate_item ::= module_or_generate_item_declaration (function_declaration)
//vparser rule name : 
//author : Codrin
//fixed by: Gabrield
module test_0250;
 (* funct = 1, test, debug *)
 function [31:0] fact;
    input in;
     fact = 32'dX;
 endfunction
endmodule
