`include "defines.v"

module b_a0(x);
// Location of source csl unit: file name = gen_uniq_rtl1.csl line number = 14
  input x;
  `include "b_a0.logic.v"
endmodule

