//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : sd_flash_lba.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module sd_flash_lba(lbdummy3,
                    lbadummy2);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 15
  input lbadummy2;
  output lbdummy3;
  `include "sd_flash_lba.logic.v"
endmodule

