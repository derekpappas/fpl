`include "defines.v"

module w0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 158
  input [1 - 1:0] ar_sa0_s10;
  v0 v0(.ar_sa0_s10(ar_sa0_s10));
  `include "w0.logic.vh"
endmodule

