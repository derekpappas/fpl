usb_tm_dispatcher.vhd
usb_tm_packetizer.vhd
usb_transaction_mgr.vhd
usb_protocol_mgr.vhd
fab.vhd
uart_mgr.vhd
RAM.vhd
jeff_uart.vhd
i2c.vhd
uart.vhd
usb_phy.vhd
fifo_regs.vhd
fab_filter.vhd
io_cell.vhd
input_cell.vhd
usb_analog_phy.vhd
output_cell.vhd
v_core.vhd
v_top.vhd
