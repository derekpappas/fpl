a.vhd
b.vhd
c.vhd
