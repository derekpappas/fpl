// Test type: always statement - loop_statement - no attribute instance
// Vparser rule name:
// Author: andreib
module alwcon16;
reg [7:0]a;
always forever a=2;
endmodule
