module testbench_output_declaration;
    output_declaration0 output_declaration_instance0();
    output_declaration1 output_declaration_instance1();
    output_declaration2 output_declaration_instance2();
    output_declaration3 output_declaration_instance3();
    output_declaration4 output_declaration_instance4();
    output_declaration5 output_declaration_instance5();
    output_declaration6 output_declaration_instance6();
    output_declaration7 output_declaration_instance7();
    output_declaration8 output_declaration_instance8();
    output_declaration9 output_declaration_instance9();
    output_declaration10 output_declaration_instance10();
    output_declaration11 output_declaration_instance11();
    output_declaration12 output_declaration_instance12();
    output_declaration13 output_declaration_instance13();
    output_declaration14 output_declaration_instance14();
    output_declaration15 output_declaration_instance15();
    output_declaration16 output_declaration_instance16();
    output_declaration17 output_declaration_instance17();
    output_declaration18 output_declaration_instance18();
    output_declaration19 output_declaration_instance19();
    output_declaration20 output_declaration_instance20();
    output_declaration21 output_declaration_instance21();
    output_declaration22 output_declaration_instance22();
    output_declaration23 output_declaration_instance23();
    output_declaration24 output_declaration_instance24();
    output_declaration25 output_declaration_instance25();
    output_declaration26 output_declaration_instance26();
    output_declaration27 output_declaration_instance27();
    output_declaration28 output_declaration_instance28();
    output_declaration29 output_declaration_instance29();
    output_declaration30 output_declaration_instance30();
    output_declaration31 output_declaration_instance31();
    output_declaration32 output_declaration_instance32();
    output_declaration33 output_declaration_instance33();
    output_declaration34 output_declaration_instance34();
    output_declaration35 output_declaration_instance35();
    output_declaration36 output_declaration_instance36();
    output_declaration37 output_declaration_instance37();
    output_declaration38 output_declaration_instance38();
    output_declaration39 output_declaration_instance39();
    output_declaration40 output_declaration_instance40();
    output_declaration41 output_declaration_instance41();
    output_declaration42 output_declaration_instance42();
    output_declaration43 output_declaration_instance43();
    output_declaration44 output_declaration_instance44();
    output_declaration45 output_declaration_instance45();
    output_declaration46 output_declaration_instance46();
    output_declaration47 output_declaration_instance47();
    output_declaration48 output_declaration_instance48();
    output_declaration49 output_declaration_instance49();
    output_declaration50 output_declaration_instance50();
    output_declaration51 output_declaration_instance51();
    output_declaration52 output_declaration_instance52();
    output_declaration53 output_declaration_instance53();
    output_declaration54 output_declaration_instance54();
    output_declaration55 output_declaration_instance55();
    output_declaration56 output_declaration_instance56();
    output_declaration57 output_declaration_instance57();
    output_declaration58 output_declaration_instance58();
    output_declaration59 output_declaration_instance59();
    output_declaration60 output_declaration_instance60();
    output_declaration61 output_declaration_instance61();
    output_declaration62 output_declaration_instance62();
    output_declaration63 output_declaration_instance63();
    output_declaration64 output_declaration_instance64();
    output_declaration65 output_declaration_instance65();
    output_declaration66 output_declaration_instance66();
    output_declaration67 output_declaration_instance67();
    output_declaration68 output_declaration_instance68();
    output_declaration69 output_declaration_instance69();
    output_declaration70 output_declaration_instance70();
    output_declaration71 output_declaration_instance71();
    output_declaration72 output_declaration_instance72();
    output_declaration73 output_declaration_instance73();
    output_declaration74 output_declaration_instance74();
    output_declaration75 output_declaration_instance75();
    output_declaration76 output_declaration_instance76();
    output_declaration77 output_declaration_instance77();
    output_declaration78 output_declaration_instance78();
    output_declaration79 output_declaration_instance79();
    output_declaration80 output_declaration_instance80();
    output_declaration81 output_declaration_instance81();
    output_declaration82 output_declaration_instance82();
    output_declaration83 output_declaration_instance83();
    output_declaration84 output_declaration_instance84();
    output_declaration85 output_declaration_instance85();
    output_declaration86 output_declaration_instance86();
    output_declaration87 output_declaration_instance87();
    output_declaration88 output_declaration_instance88();
    output_declaration89 output_declaration_instance89();
    output_declaration90 output_declaration_instance90();
    output_declaration91 output_declaration_instance91();
    output_declaration92 output_declaration_instance92();
    output_declaration93 output_declaration_instance93();
    output_declaration94 output_declaration_instance94();
    output_declaration95 output_declaration_instance95();
    output_declaration96 output_declaration_instance96();
    output_declaration97 output_declaration_instance97();
    output_declaration98 output_declaration_instance98();
    output_declaration99 output_declaration_instance99();
    output_declaration100 output_declaration_instance100();
    output_declaration101 output_declaration_instance101();
    output_declaration102 output_declaration_instance102();
    output_declaration103 output_declaration_instance103();
    output_declaration104 output_declaration_instance104();
    output_declaration105 output_declaration_instance105();
    output_declaration106 output_declaration_instance106();
    output_declaration107 output_declaration_instance107();
    output_declaration108 output_declaration_instance108();
    output_declaration109 output_declaration_instance109();
    output_declaration110 output_declaration_instance110();
    output_declaration111 output_declaration_instance111();
    output_declaration112 output_declaration_instance112();
    output_declaration113 output_declaration_instance113();
    output_declaration114 output_declaration_instance114();
    output_declaration115 output_declaration_instance115();
    output_declaration116 output_declaration_instance116();
    output_declaration117 output_declaration_instance117();
    output_declaration118 output_declaration_instance118();
    output_declaration119 output_declaration_instance119();
    output_declaration120 output_declaration_instance120();
    output_declaration121 output_declaration_instance121();
    output_declaration122 output_declaration_instance122();
    output_declaration123 output_declaration_instance123();
    output_declaration124 output_declaration_instance124();
    output_declaration125 output_declaration_instance125();
    output_declaration126 output_declaration_instance126();
    output_declaration127 output_declaration_instance127();
    output_declaration128 output_declaration_instance128();
    output_declaration129 output_declaration_instance129();
    output_declaration130 output_declaration_instance130();
    output_declaration131 output_declaration_instance131();
    output_declaration132 output_declaration_instance132();
    output_declaration133 output_declaration_instance133();
    output_declaration134 output_declaration_instance134();
    output_declaration135 output_declaration_instance135();
    output_declaration136 output_declaration_instance136();
    output_declaration137 output_declaration_instance137();
    output_declaration138 output_declaration_instance138();
    output_declaration139 output_declaration_instance139();
    output_declaration140 output_declaration_instance140();
    output_declaration141 output_declaration_instance141();
    output_declaration142 output_declaration_instance142();
    output_declaration143 output_declaration_instance143();
    output_declaration144 output_declaration_instance144();
    output_declaration145 output_declaration_instance145();
    output_declaration146 output_declaration_instance146();
    output_declaration147 output_declaration_instance147();
    output_declaration148 output_declaration_instance148();
    output_declaration149 output_declaration_instance149();
    output_declaration150 output_declaration_instance150();
    output_declaration151 output_declaration_instance151();
    output_declaration152 output_declaration_instance152();
    output_declaration153 output_declaration_instance153();
    output_declaration154 output_declaration_instance154();
    output_declaration155 output_declaration_instance155();
    output_declaration156 output_declaration_instance156();
    output_declaration157 output_declaration_instance157();
    output_declaration158 output_declaration_instance158();
    output_declaration159 output_declaration_instance159();
    output_declaration160 output_declaration_instance160();
    output_declaration161 output_declaration_instance161();
    output_declaration162 output_declaration_instance162();
    output_declaration163 output_declaration_instance163();
    output_declaration164 output_declaration_instance164();
    output_declaration165 output_declaration_instance165();
    output_declaration166 output_declaration_instance166();
    output_declaration167 output_declaration_instance167();
    output_declaration168 output_declaration_instance168();
    output_declaration169 output_declaration_instance169();
    output_declaration170 output_declaration_instance170();
    output_declaration171 output_declaration_instance171();
    output_declaration172 output_declaration_instance172();
    output_declaration173 output_declaration_instance173();
    output_declaration174 output_declaration_instance174();
    output_declaration175 output_declaration_instance175();
    output_declaration176 output_declaration_instance176();
    output_declaration177 output_declaration_instance177();
    output_declaration178 output_declaration_instance178();
    output_declaration179 output_declaration_instance179();
    output_declaration180 output_declaration_instance180();
    output_declaration181 output_declaration_instance181();
    output_declaration182 output_declaration_instance182();
    output_declaration183 output_declaration_instance183();
    output_declaration184 output_declaration_instance184();
    output_declaration185 output_declaration_instance185();
    output_declaration186 output_declaration_instance186();
    output_declaration187 output_declaration_instance187();
    output_declaration188 output_declaration_instance188();
    output_declaration189 output_declaration_instance189();
    output_declaration190 output_declaration_instance190();
    output_declaration191 output_declaration_instance191();
    output_declaration192 output_declaration_instance192();
    output_declaration193 output_declaration_instance193();
    output_declaration194 output_declaration_instance194();
    output_declaration195 output_declaration_instance195();
    output_declaration196 output_declaration_instance196();
    output_declaration197 output_declaration_instance197();
    output_declaration198 output_declaration_instance198();
    output_declaration199 output_declaration_instance199();
    output_declaration200 output_declaration_instance200();
    output_declaration201 output_declaration_instance201();
    output_declaration202 output_declaration_instance202();
    output_declaration203 output_declaration_instance203();
    output_declaration204 output_declaration_instance204();
    output_declaration205 output_declaration_instance205();
    output_declaration206 output_declaration_instance206();
    output_declaration207 output_declaration_instance207();
    output_declaration208 output_declaration_instance208();
    output_declaration209 output_declaration_instance209();
    output_declaration210 output_declaration_instance210();
    output_declaration211 output_declaration_instance211();
    output_declaration212 output_declaration_instance212();
    output_declaration213 output_declaration_instance213();
    output_declaration214 output_declaration_instance214();
    output_declaration215 output_declaration_instance215();
    output_declaration216 output_declaration_instance216();
    output_declaration217 output_declaration_instance217();
    output_declaration218 output_declaration_instance218();
    output_declaration219 output_declaration_instance219();
    output_declaration220 output_declaration_instance220();
    output_declaration221 output_declaration_instance221();
    output_declaration222 output_declaration_instance222();
    output_declaration223 output_declaration_instance223();
    output_declaration224 output_declaration_instance224();
    output_declaration225 output_declaration_instance225();
    output_declaration226 output_declaration_instance226();
    output_declaration227 output_declaration_instance227();
    output_declaration228 output_declaration_instance228();
    output_declaration229 output_declaration_instance229();
    output_declaration230 output_declaration_instance230();
    output_declaration231 output_declaration_instance231();
    output_declaration232 output_declaration_instance232();
    output_declaration233 output_declaration_instance233();
    output_declaration234 output_declaration_instance234();
    output_declaration235 output_declaration_instance235();
    output_declaration236 output_declaration_instance236();
    output_declaration237 output_declaration_instance237();
    output_declaration238 output_declaration_instance238();
    output_declaration239 output_declaration_instance239();
    output_declaration240 output_declaration_instance240();
    output_declaration241 output_declaration_instance241();
    output_declaration242 output_declaration_instance242();
    output_declaration243 output_declaration_instance243();
    output_declaration244 output_declaration_instance244();
    output_declaration245 output_declaration_instance245();
    output_declaration246 output_declaration_instance246();
    output_declaration247 output_declaration_instance247();
    output_declaration248 output_declaration_instance248();
    output_declaration249 output_declaration_instance249();
    output_declaration250 output_declaration_instance250();
    output_declaration251 output_declaration_instance251();
    output_declaration252 output_declaration_instance252();
    output_declaration253 output_declaration_instance253();
    output_declaration254 output_declaration_instance254();
    output_declaration255 output_declaration_instance255();
    output_declaration256 output_declaration_instance256();
    output_declaration257 output_declaration_instance257();
    output_declaration258 output_declaration_instance258();
    output_declaration259 output_declaration_instance259();
    output_declaration260 output_declaration_instance260();
    output_declaration261 output_declaration_instance261();
    output_declaration262 output_declaration_instance262();
    output_declaration263 output_declaration_instance263();
    output_declaration264 output_declaration_instance264();
    output_declaration265 output_declaration_instance265();
    output_declaration266 output_declaration_instance266();
    output_declaration267 output_declaration_instance267();
    output_declaration268 output_declaration_instance268();
    output_declaration269 output_declaration_instance269();
    output_declaration270 output_declaration_instance270();
    output_declaration271 output_declaration_instance271();
    output_declaration272 output_declaration_instance272();
    output_declaration273 output_declaration_instance273();
    output_declaration274 output_declaration_instance274();
    output_declaration275 output_declaration_instance275();
    output_declaration276 output_declaration_instance276();
    output_declaration277 output_declaration_instance277();
    output_declaration278 output_declaration_instance278();
    output_declaration279 output_declaration_instance279();
    output_declaration280 output_declaration_instance280();
    output_declaration281 output_declaration_instance281();
    output_declaration282 output_declaration_instance282();
    output_declaration283 output_declaration_instance283();
    output_declaration284 output_declaration_instance284();
    output_declaration285 output_declaration_instance285();
    output_declaration286 output_declaration_instance286();
    output_declaration287 output_declaration_instance287();
    output_declaration288 output_declaration_instance288();
    output_declaration289 output_declaration_instance289();
    output_declaration290 output_declaration_instance290();
    output_declaration291 output_declaration_instance291();
    output_declaration292 output_declaration_instance292();
    output_declaration293 output_declaration_instance293();
    output_declaration294 output_declaration_instance294();
    output_declaration295 output_declaration_instance295();
    output_declaration296 output_declaration_instance296();
    output_declaration297 output_declaration_instance297();
    output_declaration298 output_declaration_instance298();
    output_declaration299 output_declaration_instance299();
    output_declaration300 output_declaration_instance300();
    output_declaration301 output_declaration_instance301();
    output_declaration302 output_declaration_instance302();
    output_declaration303 output_declaration_instance303();
    output_declaration304 output_declaration_instance304();
    output_declaration305 output_declaration_instance305();
    output_declaration306 output_declaration_instance306();
    output_declaration307 output_declaration_instance307();
    output_declaration308 output_declaration_instance308();
    output_declaration309 output_declaration_instance309();
    output_declaration310 output_declaration_instance310();
    output_declaration311 output_declaration_instance311();
    output_declaration312 output_declaration_instance312();
    output_declaration313 output_declaration_instance313();
    output_declaration314 output_declaration_instance314();
    output_declaration315 output_declaration_instance315();
    output_declaration316 output_declaration_instance316();
    output_declaration317 output_declaration_instance317();
    output_declaration318 output_declaration_instance318();
    output_declaration319 output_declaration_instance319();
    output_declaration320 output_declaration_instance320();
    output_declaration321 output_declaration_instance321();
    output_declaration322 output_declaration_instance322();
    output_declaration323 output_declaration_instance323();
    output_declaration324 output_declaration_instance324();
    output_declaration325 output_declaration_instance325();
    output_declaration326 output_declaration_instance326();
    output_declaration327 output_declaration_instance327();
    output_declaration328 output_declaration_instance328();
    output_declaration329 output_declaration_instance329();
    output_declaration330 output_declaration_instance330();
    output_declaration331 output_declaration_instance331();
    output_declaration332 output_declaration_instance332();
    output_declaration333 output_declaration_instance333();
    output_declaration334 output_declaration_instance334();
    output_declaration335 output_declaration_instance335();
    output_declaration336 output_declaration_instance336();
    output_declaration337 output_declaration_instance337();
    output_declaration338 output_declaration_instance338();
    output_declaration339 output_declaration_instance339();
    output_declaration340 output_declaration_instance340();
    output_declaration341 output_declaration_instance341();
    output_declaration342 output_declaration_instance342();
    output_declaration343 output_declaration_instance343();
    output_declaration344 output_declaration_instance344();
    output_declaration345 output_declaration_instance345();
    output_declaration346 output_declaration_instance346();
    output_declaration347 output_declaration_instance347();
    output_declaration348 output_declaration_instance348();
    output_declaration349 output_declaration_instance349();
    output_declaration350 output_declaration_instance350();
    output_declaration351 output_declaration_instance351();
    output_declaration352 output_declaration_instance352();
    output_declaration353 output_declaration_instance353();
    output_declaration354 output_declaration_instance354();
    output_declaration355 output_declaration_instance355();
    output_declaration356 output_declaration_instance356();
    output_declaration357 output_declaration_instance357();
    output_declaration358 output_declaration_instance358();
    output_declaration359 output_declaration_instance359();
    output_declaration360 output_declaration_instance360();
    output_declaration361 output_declaration_instance361();
    output_declaration362 output_declaration_instance362();
    output_declaration363 output_declaration_instance363();
    output_declaration364 output_declaration_instance364();
    output_declaration365 output_declaration_instance365();
    output_declaration366 output_declaration_instance366();
    output_declaration367 output_declaration_instance367();
    output_declaration368 output_declaration_instance368();
    output_declaration369 output_declaration_instance369();
    output_declaration370 output_declaration_instance370();
    output_declaration371 output_declaration_instance371();
    output_declaration372 output_declaration_instance372();
    output_declaration373 output_declaration_instance373();
    output_declaration374 output_declaration_instance374();
    output_declaration375 output_declaration_instance375();
    output_declaration376 output_declaration_instance376();
    output_declaration377 output_declaration_instance377();
    output_declaration378 output_declaration_instance378();
    output_declaration379 output_declaration_instance379();
    output_declaration380 output_declaration_instance380();
    output_declaration381 output_declaration_instance381();
    output_declaration382 output_declaration_instance382();
    output_declaration383 output_declaration_instance383();
    output_declaration384 output_declaration_instance384();
    output_declaration385 output_declaration_instance385();
    output_declaration386 output_declaration_instance386();
    output_declaration387 output_declaration_instance387();
    output_declaration388 output_declaration_instance388();
    output_declaration389 output_declaration_instance389();
    output_declaration390 output_declaration_instance390();
    output_declaration391 output_declaration_instance391();
    output_declaration392 output_declaration_instance392();
    output_declaration393 output_declaration_instance393();
    output_declaration394 output_declaration_instance394();
    output_declaration395 output_declaration_instance395();
    output_declaration396 output_declaration_instance396();
    output_declaration397 output_declaration_instance397();
    output_declaration398 output_declaration_instance398();
    output_declaration399 output_declaration_instance399();
    output_declaration400 output_declaration_instance400();
    output_declaration401 output_declaration_instance401();
    output_declaration402 output_declaration_instance402();
    output_declaration403 output_declaration_instance403();
    output_declaration404 output_declaration_instance404();
    output_declaration405 output_declaration_instance405();
    output_declaration406 output_declaration_instance406();
    output_declaration407 output_declaration_instance407();
    output_declaration408 output_declaration_instance408();
    output_declaration409 output_declaration_instance409();
    output_declaration410 output_declaration_instance410();
    output_declaration411 output_declaration_instance411();
    output_declaration412 output_declaration_instance412();
    output_declaration413 output_declaration_instance413();
    output_declaration414 output_declaration_instance414();
    output_declaration415 output_declaration_instance415();
    output_declaration416 output_declaration_instance416();
    output_declaration417 output_declaration_instance417();
    output_declaration418 output_declaration_instance418();
    output_declaration419 output_declaration_instance419();
    output_declaration420 output_declaration_instance420();
    output_declaration421 output_declaration_instance421();
    output_declaration422 output_declaration_instance422();
    output_declaration423 output_declaration_instance423();
    output_declaration424 output_declaration_instance424();
    output_declaration425 output_declaration_instance425();
    output_declaration426 output_declaration_instance426();
    output_declaration427 output_declaration_instance427();
    output_declaration428 output_declaration_instance428();
    output_declaration429 output_declaration_instance429();
    output_declaration430 output_declaration_instance430();
    output_declaration431 output_declaration_instance431();
    output_declaration432 output_declaration_instance432();
    output_declaration433 output_declaration_instance433();
    output_declaration434 output_declaration_instance434();
    output_declaration435 output_declaration_instance435();
    output_declaration436 output_declaration_instance436();
    output_declaration437 output_declaration_instance437();
    output_declaration438 output_declaration_instance438();
    output_declaration439 output_declaration_instance439();
    output_declaration440 output_declaration_instance440();
    output_declaration441 output_declaration_instance441();
    output_declaration442 output_declaration_instance442();
    output_declaration443 output_declaration_instance443();
    output_declaration444 output_declaration_instance444();
    output_declaration445 output_declaration_instance445();
    output_declaration446 output_declaration_instance446();
    output_declaration447 output_declaration_instance447();
    output_declaration448 output_declaration_instance448();
    output_declaration449 output_declaration_instance449();
    output_declaration450 output_declaration_instance450();
    output_declaration451 output_declaration_instance451();
    output_declaration452 output_declaration_instance452();
    output_declaration453 output_declaration_instance453();
    output_declaration454 output_declaration_instance454();
    output_declaration455 output_declaration_instance455();
    output_declaration456 output_declaration_instance456();
    output_declaration457 output_declaration_instance457();
    output_declaration458 output_declaration_instance458();
    output_declaration459 output_declaration_instance459();
    output_declaration460 output_declaration_instance460();
    output_declaration461 output_declaration_instance461();
    output_declaration462 output_declaration_instance462();
    output_declaration463 output_declaration_instance463();
    output_declaration464 output_declaration_instance464();
    output_declaration465 output_declaration_instance465();
    output_declaration466 output_declaration_instance466();
    output_declaration467 output_declaration_instance467();
    output_declaration468 output_declaration_instance468();
    output_declaration469 output_declaration_instance469();
    output_declaration470 output_declaration_instance470();
    output_declaration471 output_declaration_instance471();
    output_declaration472 output_declaration_instance472();
    output_declaration473 output_declaration_instance473();
    output_declaration474 output_declaration_instance474();
    output_declaration475 output_declaration_instance475();
    output_declaration476 output_declaration_instance476();
    output_declaration477 output_declaration_instance477();
    output_declaration478 output_declaration_instance478();
    output_declaration479 output_declaration_instance479();
    output_declaration480 output_declaration_instance480();
    output_declaration481 output_declaration_instance481();
    output_declaration482 output_declaration_instance482();
    output_declaration483 output_declaration_instance483();
    output_declaration484 output_declaration_instance484();
    output_declaration485 output_declaration_instance485();
    output_declaration486 output_declaration_instance486();
    output_declaration487 output_declaration_instance487();
    output_declaration488 output_declaration_instance488();
    output_declaration489 output_declaration_instance489();
    output_declaration490 output_declaration_instance490();
    output_declaration491 output_declaration_instance491();
    output_declaration492 output_declaration_instance492();
    output_declaration493 output_declaration_instance493();
    output_declaration494 output_declaration_instance494();
    output_declaration495 output_declaration_instance495();
    output_declaration496 output_declaration_instance496();
    output_declaration497 output_declaration_instance497();
    output_declaration498 output_declaration_instance498();
    output_declaration499 output_declaration_instance499();
    output_declaration500 output_declaration_instance500();
    output_declaration501 output_declaration_instance501();
    output_declaration502 output_declaration_instance502();
    output_declaration503 output_declaration_instance503();
    output_declaration504 output_declaration_instance504();
    output_declaration505 output_declaration_instance505();
    output_declaration506 output_declaration_instance506();
    output_declaration507 output_declaration_instance507();
    output_declaration508 output_declaration_instance508();
    output_declaration509 output_declaration_instance509();
    output_declaration510 output_declaration_instance510();
    output_declaration511 output_declaration_instance511();
    output_declaration512 output_declaration_instance512();
    output_declaration513 output_declaration_instance513();
    output_declaration514 output_declaration_instance514();
    output_declaration515 output_declaration_instance515();
    output_declaration516 output_declaration_instance516();
    output_declaration517 output_declaration_instance517();
    output_declaration518 output_declaration_instance518();
    output_declaration519 output_declaration_instance519();
    output_declaration520 output_declaration_instance520();
    output_declaration521 output_declaration_instance521();
    output_declaration522 output_declaration_instance522();
    output_declaration523 output_declaration_instance523();
    output_declaration524 output_declaration_instance524();
    output_declaration525 output_declaration_instance525();
    output_declaration526 output_declaration_instance526();
    output_declaration527 output_declaration_instance527();
    output_declaration528 output_declaration_instance528();
    output_declaration529 output_declaration_instance529();
    output_declaration530 output_declaration_instance530();
    output_declaration531 output_declaration_instance531();
    output_declaration532 output_declaration_instance532();
    output_declaration533 output_declaration_instance533();
    output_declaration534 output_declaration_instance534();
    output_declaration535 output_declaration_instance535();
    output_declaration536 output_declaration_instance536();
    output_declaration537 output_declaration_instance537();
    output_declaration538 output_declaration_instance538();
    output_declaration539 output_declaration_instance539();
    output_declaration540 output_declaration_instance540();
    output_declaration541 output_declaration_instance541();
    output_declaration542 output_declaration_instance542();
    output_declaration543 output_declaration_instance543();
    output_declaration544 output_declaration_instance544();
    output_declaration545 output_declaration_instance545();
    output_declaration546 output_declaration_instance546();
    output_declaration547 output_declaration_instance547();
    output_declaration548 output_declaration_instance548();
    output_declaration549 output_declaration_instance549();
    output_declaration550 output_declaration_instance550();
    output_declaration551 output_declaration_instance551();
    output_declaration552 output_declaration_instance552();
    output_declaration553 output_declaration_instance553();
    output_declaration554 output_declaration_instance554();
    output_declaration555 output_declaration_instance555();
    output_declaration556 output_declaration_instance556();
    output_declaration557 output_declaration_instance557();
    output_declaration558 output_declaration_instance558();
    output_declaration559 output_declaration_instance559();
    output_declaration560 output_declaration_instance560();
    output_declaration561 output_declaration_instance561();
    output_declaration562 output_declaration_instance562();
    output_declaration563 output_declaration_instance563();
    output_declaration564 output_declaration_instance564();
    output_declaration565 output_declaration_instance565();
    output_declaration566 output_declaration_instance566();
    output_declaration567 output_declaration_instance567();
    output_declaration568 output_declaration_instance568();
    output_declaration569 output_declaration_instance569();
    output_declaration570 output_declaration_instance570();
    output_declaration571 output_declaration_instance571();
    output_declaration572 output_declaration_instance572();
    output_declaration573 output_declaration_instance573();
    output_declaration574 output_declaration_instance574();
    output_declaration575 output_declaration_instance575();
    output_declaration576 output_declaration_instance576();
    output_declaration577 output_declaration_instance577();
    output_declaration578 output_declaration_instance578();
    output_declaration579 output_declaration_instance579();
    output_declaration580 output_declaration_instance580();
    output_declaration581 output_declaration_instance581();
    output_declaration582 output_declaration_instance582();
    output_declaration583 output_declaration_instance583();
    output_declaration584 output_declaration_instance584();
    output_declaration585 output_declaration_instance585();
    output_declaration586 output_declaration_instance586();
    output_declaration587 output_declaration_instance587();
    output_declaration588 output_declaration_instance588();
    output_declaration589 output_declaration_instance589();
    output_declaration590 output_declaration_instance590();
    output_declaration591 output_declaration_instance591();
    output_declaration592 output_declaration_instance592();
    output_declaration593 output_declaration_instance593();
    output_declaration594 output_declaration_instance594();
    output_declaration595 output_declaration_instance595();
    output_declaration596 output_declaration_instance596();
    output_declaration597 output_declaration_instance597();
    output_declaration598 output_declaration_instance598();
    output_declaration599 output_declaration_instance599();
    output_declaration600 output_declaration_instance600();
    output_declaration601 output_declaration_instance601();
    output_declaration602 output_declaration_instance602();
    output_declaration603 output_declaration_instance603();
    output_declaration604 output_declaration_instance604();
    output_declaration605 output_declaration_instance605();
    output_declaration606 output_declaration_instance606();
    output_declaration607 output_declaration_instance607();
    output_declaration608 output_declaration_instance608();
    output_declaration609 output_declaration_instance609();
    output_declaration610 output_declaration_instance610();
    output_declaration611 output_declaration_instance611();
    output_declaration612 output_declaration_instance612();
    output_declaration613 output_declaration_instance613();
    output_declaration614 output_declaration_instance614();
    output_declaration615 output_declaration_instance615();
    output_declaration616 output_declaration_instance616();
    output_declaration617 output_declaration_instance617();
    output_declaration618 output_declaration_instance618();
    output_declaration619 output_declaration_instance619();
    output_declaration620 output_declaration_instance620();
    output_declaration621 output_declaration_instance621();
    output_declaration622 output_declaration_instance622();
    output_declaration623 output_declaration_instance623();
    output_declaration624 output_declaration_instance624();
    output_declaration625 output_declaration_instance625();
    output_declaration626 output_declaration_instance626();
    output_declaration627 output_declaration_instance627();
    output_declaration628 output_declaration_instance628();
    output_declaration629 output_declaration_instance629();
    output_declaration630 output_declaration_instance630();
    output_declaration631 output_declaration_instance631();
    output_declaration632 output_declaration_instance632();
    output_declaration633 output_declaration_instance633();
    output_declaration634 output_declaration_instance634();
    output_declaration635 output_declaration_instance635();
    output_declaration636 output_declaration_instance636();
    output_declaration637 output_declaration_instance637();
    output_declaration638 output_declaration_instance638();
    output_declaration639 output_declaration_instance639();
    output_declaration640 output_declaration_instance640();
    output_declaration641 output_declaration_instance641();
    output_declaration642 output_declaration_instance642();
    output_declaration643 output_declaration_instance643();
    output_declaration644 output_declaration_instance644();
    output_declaration645 output_declaration_instance645();
    output_declaration646 output_declaration_instance646();
    output_declaration647 output_declaration_instance647();
    output_declaration648 output_declaration_instance648();
    output_declaration649 output_declaration_instance649();
    output_declaration650 output_declaration_instance650();
    output_declaration651 output_declaration_instance651();
    output_declaration652 output_declaration_instance652();
    output_declaration653 output_declaration_instance653();
    output_declaration654 output_declaration_instance654();
    output_declaration655 output_declaration_instance655();
    output_declaration656 output_declaration_instance656();
    output_declaration657 output_declaration_instance657();
    output_declaration658 output_declaration_instance658();
    output_declaration659 output_declaration_instance659();
    output_declaration660 output_declaration_instance660();
    output_declaration661 output_declaration_instance661();
    output_declaration662 output_declaration_instance662();
    output_declaration663 output_declaration_instance663();
    output_declaration664 output_declaration_instance664();
    output_declaration665 output_declaration_instance665();
    output_declaration666 output_declaration_instance666();
    output_declaration667 output_declaration_instance667();
    output_declaration668 output_declaration_instance668();
    output_declaration669 output_declaration_instance669();
    output_declaration670 output_declaration_instance670();
    output_declaration671 output_declaration_instance671();
    output_declaration672 output_declaration_instance672();
    output_declaration673 output_declaration_instance673();
    output_declaration674 output_declaration_instance674();
    output_declaration675 output_declaration_instance675();
    output_declaration676 output_declaration_instance676();
    output_declaration677 output_declaration_instance677();
    output_declaration678 output_declaration_instance678();
    output_declaration679 output_declaration_instance679();
    output_declaration680 output_declaration_instance680();
    output_declaration681 output_declaration_instance681();
    output_declaration682 output_declaration_instance682();
    output_declaration683 output_declaration_instance683();
    output_declaration684 output_declaration_instance684();
    output_declaration685 output_declaration_instance685();
    output_declaration686 output_declaration_instance686();
    output_declaration687 output_declaration_instance687();
    output_declaration688 output_declaration_instance688();
    output_declaration689 output_declaration_instance689();
    output_declaration690 output_declaration_instance690();
    output_declaration691 output_declaration_instance691();
    output_declaration692 output_declaration_instance692();
    output_declaration693 output_declaration_instance693();
    output_declaration694 output_declaration_instance694();
    output_declaration695 output_declaration_instance695();
    output_declaration696 output_declaration_instance696();
    output_declaration697 output_declaration_instance697();
    output_declaration698 output_declaration_instance698();
    output_declaration699 output_declaration_instance699();
    output_declaration700 output_declaration_instance700();
    output_declaration701 output_declaration_instance701();
    output_declaration702 output_declaration_instance702();
    output_declaration703 output_declaration_instance703();
    output_declaration704 output_declaration_instance704();
    output_declaration705 output_declaration_instance705();
    output_declaration706 output_declaration_instance706();
    output_declaration707 output_declaration_instance707();
    output_declaration708 output_declaration_instance708();
    output_declaration709 output_declaration_instance709();
    output_declaration710 output_declaration_instance710();
    output_declaration711 output_declaration_instance711();
    output_declaration712 output_declaration_instance712();
    output_declaration713 output_declaration_instance713();
    output_declaration714 output_declaration_instance714();
    output_declaration715 output_declaration_instance715();
    output_declaration716 output_declaration_instance716();
    output_declaration717 output_declaration_instance717();
    output_declaration718 output_declaration_instance718();
    output_declaration719 output_declaration_instance719();
    output_declaration720 output_declaration_instance720();
    output_declaration721 output_declaration_instance721();
    output_declaration722 output_declaration_instance722();
    output_declaration723 output_declaration_instance723();
    output_declaration724 output_declaration_instance724();
    output_declaration725 output_declaration_instance725();
    output_declaration726 output_declaration_instance726();
    output_declaration727 output_declaration_instance727();
    output_declaration728 output_declaration_instance728();
    output_declaration729 output_declaration_instance729();
    output_declaration730 output_declaration_instance730();
    output_declaration731 output_declaration_instance731();
    output_declaration732 output_declaration_instance732();
    output_declaration733 output_declaration_instance733();
    output_declaration734 output_declaration_instance734();
    output_declaration735 output_declaration_instance735();
    output_declaration736 output_declaration_instance736();
    output_declaration737 output_declaration_instance737();
    output_declaration738 output_declaration_instance738();
    output_declaration739 output_declaration_instance739();
    output_declaration740 output_declaration_instance740();
    output_declaration741 output_declaration_instance741();
    output_declaration742 output_declaration_instance742();
    output_declaration743 output_declaration_instance743();
    output_declaration744 output_declaration_instance744();
    output_declaration745 output_declaration_instance745();
    output_declaration746 output_declaration_instance746();
    output_declaration747 output_declaration_instance747();
    output_declaration748 output_declaration_instance748();
    output_declaration749 output_declaration_instance749();
    output_declaration750 output_declaration_instance750();
    output_declaration751 output_declaration_instance751();
    output_declaration752 output_declaration_instance752();
    output_declaration753 output_declaration_instance753();
    output_declaration754 output_declaration_instance754();
    output_declaration755 output_declaration_instance755();
    output_declaration756 output_declaration_instance756();
    output_declaration757 output_declaration_instance757();
    output_declaration758 output_declaration_instance758();
    output_declaration759 output_declaration_instance759();
    output_declaration760 output_declaration_instance760();
    output_declaration761 output_declaration_instance761();
    output_declaration762 output_declaration_instance762();
    output_declaration763 output_declaration_instance763();
    output_declaration764 output_declaration_instance764();
    output_declaration765 output_declaration_instance765();
    output_declaration766 output_declaration_instance766();
    output_declaration767 output_declaration_instance767();
    output_declaration768 output_declaration_instance768();
    output_declaration769 output_declaration_instance769();
    output_declaration770 output_declaration_instance770();
    output_declaration771 output_declaration_instance771();
    output_declaration772 output_declaration_instance772();
    output_declaration773 output_declaration_instance773();
    output_declaration774 output_declaration_instance774();
    output_declaration775 output_declaration_instance775();
    output_declaration776 output_declaration_instance776();
    output_declaration777 output_declaration_instance777();
    output_declaration778 output_declaration_instance778();
    output_declaration779 output_declaration_instance779();
    output_declaration780 output_declaration_instance780();
    output_declaration781 output_declaration_instance781();
    output_declaration782 output_declaration_instance782();
    output_declaration783 output_declaration_instance783();
    output_declaration784 output_declaration_instance784();
    output_declaration785 output_declaration_instance785();
    output_declaration786 output_declaration_instance786();
    output_declaration787 output_declaration_instance787();
    output_declaration788 output_declaration_instance788();
    output_declaration789 output_declaration_instance789();
    output_declaration790 output_declaration_instance790();
    output_declaration791 output_declaration_instance791();
    output_declaration792 output_declaration_instance792();
    output_declaration793 output_declaration_instance793();
    output_declaration794 output_declaration_instance794();
    output_declaration795 output_declaration_instance795();
    output_declaration796 output_declaration_instance796();
    output_declaration797 output_declaration_instance797();
    output_declaration798 output_declaration_instance798();
    output_declaration799 output_declaration_instance799();
    output_declaration800 output_declaration_instance800();
    output_declaration801 output_declaration_instance801();
    output_declaration802 output_declaration_instance802();
    output_declaration803 output_declaration_instance803();
    output_declaration804 output_declaration_instance804();
    output_declaration805 output_declaration_instance805();
    output_declaration806 output_declaration_instance806();
    output_declaration807 output_declaration_instance807();
    output_declaration808 output_declaration_instance808();
    output_declaration809 output_declaration_instance809();
    output_declaration810 output_declaration_instance810();
    output_declaration811 output_declaration_instance811();
    output_declaration812 output_declaration_instance812();
    output_declaration813 output_declaration_instance813();
    output_declaration814 output_declaration_instance814();
    output_declaration815 output_declaration_instance815();
    output_declaration816 output_declaration_instance816();
    output_declaration817 output_declaration_instance817();
    output_declaration818 output_declaration_instance818();
    output_declaration819 output_declaration_instance819();
    output_declaration820 output_declaration_instance820();
    output_declaration821 output_declaration_instance821();
    output_declaration822 output_declaration_instance822();
    output_declaration823 output_declaration_instance823();
    output_declaration824 output_declaration_instance824();
    output_declaration825 output_declaration_instance825();
    output_declaration826 output_declaration_instance826();
    output_declaration827 output_declaration_instance827();
    output_declaration828 output_declaration_instance828();
    output_declaration829 output_declaration_instance829();
    output_declaration830 output_declaration_instance830();
    output_declaration831 output_declaration_instance831();
    output_declaration832 output_declaration_instance832();
    output_declaration833 output_declaration_instance833();
    output_declaration834 output_declaration_instance834();
    output_declaration835 output_declaration_instance835();
    output_declaration836 output_declaration_instance836();
    output_declaration837 output_declaration_instance837();
    output_declaration838 output_declaration_instance838();
    output_declaration839 output_declaration_instance839();
    output_declaration840 output_declaration_instance840();
    output_declaration841 output_declaration_instance841();
    output_declaration842 output_declaration_instance842();
    output_declaration843 output_declaration_instance843();
    output_declaration844 output_declaration_instance844();
    output_declaration845 output_declaration_instance845();
    output_declaration846 output_declaration_instance846();
    output_declaration847 output_declaration_instance847();
    output_declaration848 output_declaration_instance848();
    output_declaration849 output_declaration_instance849();
    output_declaration850 output_declaration_instance850();
    output_declaration851 output_declaration_instance851();
    output_declaration852 output_declaration_instance852();
    output_declaration853 output_declaration_instance853();
    output_declaration854 output_declaration_instance854();
    output_declaration855 output_declaration_instance855();
    output_declaration856 output_declaration_instance856();
    output_declaration857 output_declaration_instance857();
    output_declaration858 output_declaration_instance858();
    output_declaration859 output_declaration_instance859();
    output_declaration860 output_declaration_instance860();
    output_declaration861 output_declaration_instance861();
    output_declaration862 output_declaration_instance862();
    output_declaration863 output_declaration_instance863();
    output_declaration864 output_declaration_instance864();
    output_declaration865 output_declaration_instance865();
    output_declaration866 output_declaration_instance866();
    output_declaration867 output_declaration_instance867();
    output_declaration868 output_declaration_instance868();
    output_declaration869 output_declaration_instance869();
    output_declaration870 output_declaration_instance870();
    output_declaration871 output_declaration_instance871();
    output_declaration872 output_declaration_instance872();
    output_declaration873 output_declaration_instance873();
    output_declaration874 output_declaration_instance874();
    output_declaration875 output_declaration_instance875();
    output_declaration876 output_declaration_instance876();
    output_declaration877 output_declaration_instance877();
    output_declaration878 output_declaration_instance878();
    output_declaration879 output_declaration_instance879();
    output_declaration880 output_declaration_instance880();
    output_declaration881 output_declaration_instance881();
    output_declaration882 output_declaration_instance882();
    output_declaration883 output_declaration_instance883();
    output_declaration884 output_declaration_instance884();
    output_declaration885 output_declaration_instance885();
    output_declaration886 output_declaration_instance886();
    output_declaration887 output_declaration_instance887();
    output_declaration888 output_declaration_instance888();
    output_declaration889 output_declaration_instance889();
    output_declaration890 output_declaration_instance890();
    output_declaration891 output_declaration_instance891();
    output_declaration892 output_declaration_instance892();
    output_declaration893 output_declaration_instance893();
    output_declaration894 output_declaration_instance894();
    output_declaration895 output_declaration_instance895();
    output_declaration896 output_declaration_instance896();
    output_declaration897 output_declaration_instance897();
    output_declaration898 output_declaration_instance898();
    output_declaration899 output_declaration_instance899();
    output_declaration900 output_declaration_instance900();
    output_declaration901 output_declaration_instance901();
    output_declaration902 output_declaration_instance902();
    output_declaration903 output_declaration_instance903();
    output_declaration904 output_declaration_instance904();
    output_declaration905 output_declaration_instance905();
    output_declaration906 output_declaration_instance906();
    output_declaration907 output_declaration_instance907();
    output_declaration908 output_declaration_instance908();
    output_declaration909 output_declaration_instance909();
    output_declaration910 output_declaration_instance910();
    output_declaration911 output_declaration_instance911();
    output_declaration912 output_declaration_instance912();
    output_declaration913 output_declaration_instance913();
    output_declaration914 output_declaration_instance914();
    output_declaration915 output_declaration_instance915();
    output_declaration916 output_declaration_instance916();
    output_declaration917 output_declaration_instance917();
    output_declaration918 output_declaration_instance918();
    output_declaration919 output_declaration_instance919();
    output_declaration920 output_declaration_instance920();
    output_declaration921 output_declaration_instance921();
    output_declaration922 output_declaration_instance922();
    output_declaration923 output_declaration_instance923();
    output_declaration924 output_declaration_instance924();
    output_declaration925 output_declaration_instance925();
    output_declaration926 output_declaration_instance926();
    output_declaration927 output_declaration_instance927();
    output_declaration928 output_declaration_instance928();
    output_declaration929 output_declaration_instance929();
    output_declaration930 output_declaration_instance930();
    output_declaration931 output_declaration_instance931();
    output_declaration932 output_declaration_instance932();
    output_declaration933 output_declaration_instance933();
    output_declaration934 output_declaration_instance934();
    output_declaration935 output_declaration_instance935();
    output_declaration936 output_declaration_instance936();
    output_declaration937 output_declaration_instance937();
    output_declaration938 output_declaration_instance938();
    output_declaration939 output_declaration_instance939();
    output_declaration940 output_declaration_instance940();
    output_declaration941 output_declaration_instance941();
    output_declaration942 output_declaration_instance942();
    output_declaration943 output_declaration_instance943();
    output_declaration944 output_declaration_instance944();
    output_declaration945 output_declaration_instance945();
    output_declaration946 output_declaration_instance946();
    output_declaration947 output_declaration_instance947();
    output_declaration948 output_declaration_instance948();
    output_declaration949 output_declaration_instance949();
    output_declaration950 output_declaration_instance950();
    output_declaration951 output_declaration_instance951();
    output_declaration952 output_declaration_instance952();
    output_declaration953 output_declaration_instance953();
    output_declaration954 output_declaration_instance954();
    output_declaration955 output_declaration_instance955();
    output_declaration956 output_declaration_instance956();
    output_declaration957 output_declaration_instance957();
    output_declaration958 output_declaration_instance958();
    output_declaration959 output_declaration_instance959();
    output_declaration960 output_declaration_instance960();
    output_declaration961 output_declaration_instance961();
    output_declaration962 output_declaration_instance962();
    output_declaration963 output_declaration_instance963();
    output_declaration964 output_declaration_instance964();
    output_declaration965 output_declaration_instance965();
    output_declaration966 output_declaration_instance966();
    output_declaration967 output_declaration_instance967();
    output_declaration968 output_declaration_instance968();
    output_declaration969 output_declaration_instance969();
    output_declaration970 output_declaration_instance970();
    output_declaration971 output_declaration_instance971();
    output_declaration972 output_declaration_instance972();
    output_declaration973 output_declaration_instance973();
    output_declaration974 output_declaration_instance974();
    output_declaration975 output_declaration_instance975();
    output_declaration976 output_declaration_instance976();
    output_declaration977 output_declaration_instance977();
    output_declaration978 output_declaration_instance978();
    output_declaration979 output_declaration_instance979();
    output_declaration980 output_declaration_instance980();
    output_declaration981 output_declaration_instance981();
    output_declaration982 output_declaration_instance982();
    output_declaration983 output_declaration_instance983();
    output_declaration984 output_declaration_instance984();
    output_declaration985 output_declaration_instance985();
    output_declaration986 output_declaration_instance986();
    output_declaration987 output_declaration_instance987();
    output_declaration988 output_declaration_instance988();
    output_declaration989 output_declaration_instance989();
    output_declaration990 output_declaration_instance990();
    output_declaration991 output_declaration_instance991();
    output_declaration992 output_declaration_instance992();
    output_declaration993 output_declaration_instance993();
    output_declaration994 output_declaration_instance994();
    output_declaration995 output_declaration_instance995();
    output_declaration996 output_declaration_instance996();
    output_declaration997 output_declaration_instance997();
    output_declaration998 output_declaration_instance998();
    output_declaration999 output_declaration_instance999();
    output_declaration1000 output_declaration_instance1000();
    output_declaration1001 output_declaration_instance1001();
    output_declaration1002 output_declaration_instance1002();
    output_declaration1003 output_declaration_instance1003();
    output_declaration1004 output_declaration_instance1004();
    output_declaration1005 output_declaration_instance1005();
    output_declaration1006 output_declaration_instance1006();
    output_declaration1007 output_declaration_instance1007();
    output_declaration1008 output_declaration_instance1008();
    output_declaration1009 output_declaration_instance1009();
    output_declaration1010 output_declaration_instance1010();
    output_declaration1011 output_declaration_instance1011();
    output_declaration1012 output_declaration_instance1012();
    output_declaration1013 output_declaration_instance1013();
    output_declaration1014 output_declaration_instance1014();
    output_declaration1015 output_declaration_instance1015();
    output_declaration1016 output_declaration_instance1016();
    output_declaration1017 output_declaration_instance1017();
    output_declaration1018 output_declaration_instance1018();
    output_declaration1019 output_declaration_instance1019();
    output_declaration1020 output_declaration_instance1020();
    output_declaration1021 output_declaration_instance1021();
    output_declaration1022 output_declaration_instance1022();
    output_declaration1023 output_declaration_instance1023();
    output_declaration1024 output_declaration_instance1024();
    output_declaration1025 output_declaration_instance1025();
    output_declaration1026 output_declaration_instance1026();
    output_declaration1027 output_declaration_instance1027();
    output_declaration1028 output_declaration_instance1028();
    output_declaration1029 output_declaration_instance1029();
    output_declaration1030 output_declaration_instance1030();
    output_declaration1031 output_declaration_instance1031();
    output_declaration1032 output_declaration_instance1032();
    output_declaration1033 output_declaration_instance1033();
    output_declaration1034 output_declaration_instance1034();
    output_declaration1035 output_declaration_instance1035();
    output_declaration1036 output_declaration_instance1036();
    output_declaration1037 output_declaration_instance1037();
    output_declaration1038 output_declaration_instance1038();
    output_declaration1039 output_declaration_instance1039();
    output_declaration1040 output_declaration_instance1040();
    output_declaration1041 output_declaration_instance1041();
    output_declaration1042 output_declaration_instance1042();
    output_declaration1043 output_declaration_instance1043();
    output_declaration1044 output_declaration_instance1044();
    output_declaration1045 output_declaration_instance1045();
    output_declaration1046 output_declaration_instance1046();
    output_declaration1047 output_declaration_instance1047();
    output_declaration1048 output_declaration_instance1048();
    output_declaration1049 output_declaration_instance1049();
    output_declaration1050 output_declaration_instance1050();
    output_declaration1051 output_declaration_instance1051();
    output_declaration1052 output_declaration_instance1052();
    output_declaration1053 output_declaration_instance1053();
    output_declaration1054 output_declaration_instance1054();
    output_declaration1055 output_declaration_instance1055();
    output_declaration1056 output_declaration_instance1056();
    output_declaration1057 output_declaration_instance1057();
    output_declaration1058 output_declaration_instance1058();
    output_declaration1059 output_declaration_instance1059();
    output_declaration1060 output_declaration_instance1060();
    output_declaration1061 output_declaration_instance1061();
    output_declaration1062 output_declaration_instance1062();
    output_declaration1063 output_declaration_instance1063();
    output_declaration1064 output_declaration_instance1064();
    output_declaration1065 output_declaration_instance1065();
    output_declaration1066 output_declaration_instance1066();
    output_declaration1067 output_declaration_instance1067();
    output_declaration1068 output_declaration_instance1068();
    output_declaration1069 output_declaration_instance1069();
    output_declaration1070 output_declaration_instance1070();
    output_declaration1071 output_declaration_instance1071();
    output_declaration1072 output_declaration_instance1072();
    output_declaration1073 output_declaration_instance1073();
    output_declaration1074 output_declaration_instance1074();
    output_declaration1075 output_declaration_instance1075();
    output_declaration1076 output_declaration_instance1076();
    output_declaration1077 output_declaration_instance1077();
    output_declaration1078 output_declaration_instance1078();
    output_declaration1079 output_declaration_instance1079();
    output_declaration1080 output_declaration_instance1080();
    output_declaration1081 output_declaration_instance1081();
    output_declaration1082 output_declaration_instance1082();
    output_declaration1083 output_declaration_instance1083();
    output_declaration1084 output_declaration_instance1084();
    output_declaration1085 output_declaration_instance1085();
    output_declaration1086 output_declaration_instance1086();
    output_declaration1087 output_declaration_instance1087();
    output_declaration1088 output_declaration_instance1088();
    output_declaration1089 output_declaration_instance1089();
    output_declaration1090 output_declaration_instance1090();
    output_declaration1091 output_declaration_instance1091();
    output_declaration1092 output_declaration_instance1092();
    output_declaration1093 output_declaration_instance1093();
    output_declaration1094 output_declaration_instance1094();
    output_declaration1095 output_declaration_instance1095();
    output_declaration1096 output_declaration_instance1096();
    output_declaration1097 output_declaration_instance1097();
    output_declaration1098 output_declaration_instance1098();
    output_declaration1099 output_declaration_instance1099();
    output_declaration1100 output_declaration_instance1100();
    output_declaration1101 output_declaration_instance1101();
    output_declaration1102 output_declaration_instance1102();
    output_declaration1103 output_declaration_instance1103();
    output_declaration1104 output_declaration_instance1104();
    output_declaration1105 output_declaration_instance1105();
    output_declaration1106 output_declaration_instance1106();
    output_declaration1107 output_declaration_instance1107();
    output_declaration1108 output_declaration_instance1108();
    output_declaration1109 output_declaration_instance1109();
    output_declaration1110 output_declaration_instance1110();
    output_declaration1111 output_declaration_instance1111();
    output_declaration1112 output_declaration_instance1112();
    output_declaration1113 output_declaration_instance1113();
    output_declaration1114 output_declaration_instance1114();
    output_declaration1115 output_declaration_instance1115();
    output_declaration1116 output_declaration_instance1116();
    output_declaration1117 output_declaration_instance1117();
    output_declaration1118 output_declaration_instance1118();
    output_declaration1119 output_declaration_instance1119();
    output_declaration1120 output_declaration_instance1120();
    output_declaration1121 output_declaration_instance1121();
    output_declaration1122 output_declaration_instance1122();
    output_declaration1123 output_declaration_instance1123();
    output_declaration1124 output_declaration_instance1124();
    output_declaration1125 output_declaration_instance1125();
    output_declaration1126 output_declaration_instance1126();
    output_declaration1127 output_declaration_instance1127();
    output_declaration1128 output_declaration_instance1128();
    output_declaration1129 output_declaration_instance1129();
    output_declaration1130 output_declaration_instance1130();
    output_declaration1131 output_declaration_instance1131();
    output_declaration1132 output_declaration_instance1132();
    output_declaration1133 output_declaration_instance1133();
    output_declaration1134 output_declaration_instance1134();
    output_declaration1135 output_declaration_instance1135();
    output_declaration1136 output_declaration_instance1136();
    output_declaration1137 output_declaration_instance1137();
    output_declaration1138 output_declaration_instance1138();
    output_declaration1139 output_declaration_instance1139();
    output_declaration1140 output_declaration_instance1140();
    output_declaration1141 output_declaration_instance1141();
    output_declaration1142 output_declaration_instance1142();
    output_declaration1143 output_declaration_instance1143();
    output_declaration1144 output_declaration_instance1144();
    output_declaration1145 output_declaration_instance1145();
    output_declaration1146 output_declaration_instance1146();
    output_declaration1147 output_declaration_instance1147();
    output_declaration1148 output_declaration_instance1148();
    output_declaration1149 output_declaration_instance1149();
    output_declaration1150 output_declaration_instance1150();
    output_declaration1151 output_declaration_instance1151();
    output_declaration1152 output_declaration_instance1152();
    output_declaration1153 output_declaration_instance1153();
    output_declaration1154 output_declaration_instance1154();
    output_declaration1155 output_declaration_instance1155();
    output_declaration1156 output_declaration_instance1156();
    output_declaration1157 output_declaration_instance1157();
    output_declaration1158 output_declaration_instance1158();
    output_declaration1159 output_declaration_instance1159();
    output_declaration1160 output_declaration_instance1160();
    output_declaration1161 output_declaration_instance1161();
    output_declaration1162 output_declaration_instance1162();
    output_declaration1163 output_declaration_instance1163();
    output_declaration1164 output_declaration_instance1164();
    output_declaration1165 output_declaration_instance1165();
    output_declaration1166 output_declaration_instance1166();
    output_declaration1167 output_declaration_instance1167();
    output_declaration1168 output_declaration_instance1168();
    output_declaration1169 output_declaration_instance1169();
    output_declaration1170 output_declaration_instance1170();
    output_declaration1171 output_declaration_instance1171();
    output_declaration1172 output_declaration_instance1172();
    output_declaration1173 output_declaration_instance1173();
    output_declaration1174 output_declaration_instance1174();
    output_declaration1175 output_declaration_instance1175();
    output_declaration1176 output_declaration_instance1176();
    output_declaration1177 output_declaration_instance1177();
    output_declaration1178 output_declaration_instance1178();
    output_declaration1179 output_declaration_instance1179();
    output_declaration1180 output_declaration_instance1180();
    output_declaration1181 output_declaration_instance1181();
    output_declaration1182 output_declaration_instance1182();
    output_declaration1183 output_declaration_instance1183();
    output_declaration1184 output_declaration_instance1184();
    output_declaration1185 output_declaration_instance1185();
    output_declaration1186 output_declaration_instance1186();
    output_declaration1187 output_declaration_instance1187();
    output_declaration1188 output_declaration_instance1188();
    output_declaration1189 output_declaration_instance1189();
    output_declaration1190 output_declaration_instance1190();
    output_declaration1191 output_declaration_instance1191();
    output_declaration1192 output_declaration_instance1192();
    output_declaration1193 output_declaration_instance1193();
    output_declaration1194 output_declaration_instance1194();
    output_declaration1195 output_declaration_instance1195();
    output_declaration1196 output_declaration_instance1196();
    output_declaration1197 output_declaration_instance1197();
    output_declaration1198 output_declaration_instance1198();
    output_declaration1199 output_declaration_instance1199();
    output_declaration1200 output_declaration_instance1200();
    output_declaration1201 output_declaration_instance1201();
    output_declaration1202 output_declaration_instance1202();
    output_declaration1203 output_declaration_instance1203();
    output_declaration1204 output_declaration_instance1204();
    output_declaration1205 output_declaration_instance1205();
    output_declaration1206 output_declaration_instance1206();
    output_declaration1207 output_declaration_instance1207();
    output_declaration1208 output_declaration_instance1208();
    output_declaration1209 output_declaration_instance1209();
    output_declaration1210 output_declaration_instance1210();
    output_declaration1211 output_declaration_instance1211();
    output_declaration1212 output_declaration_instance1212();
    output_declaration1213 output_declaration_instance1213();
    output_declaration1214 output_declaration_instance1214();
    output_declaration1215 output_declaration_instance1215();
    output_declaration1216 output_declaration_instance1216();
    output_declaration1217 output_declaration_instance1217();
    output_declaration1218 output_declaration_instance1218();
    output_declaration1219 output_declaration_instance1219();
    output_declaration1220 output_declaration_instance1220();
    output_declaration1221 output_declaration_instance1221();
    output_declaration1222 output_declaration_instance1222();
    output_declaration1223 output_declaration_instance1223();
    output_declaration1224 output_declaration_instance1224();
    output_declaration1225 output_declaration_instance1225();
    output_declaration1226 output_declaration_instance1226();
    output_declaration1227 output_declaration_instance1227();
    output_declaration1228 output_declaration_instance1228();
    output_declaration1229 output_declaration_instance1229();
    output_declaration1230 output_declaration_instance1230();
    output_declaration1231 output_declaration_instance1231();
    output_declaration1232 output_declaration_instance1232();
    output_declaration1233 output_declaration_instance1233();
    output_declaration1234 output_declaration_instance1234();
    output_declaration1235 output_declaration_instance1235();
    output_declaration1236 output_declaration_instance1236();
    output_declaration1237 output_declaration_instance1237();
    output_declaration1238 output_declaration_instance1238();
    output_declaration1239 output_declaration_instance1239();
    output_declaration1240 output_declaration_instance1240();
    output_declaration1241 output_declaration_instance1241();
    output_declaration1242 output_declaration_instance1242();
    output_declaration1243 output_declaration_instance1243();
    output_declaration1244 output_declaration_instance1244();
    output_declaration1245 output_declaration_instance1245();
    output_declaration1246 output_declaration_instance1246();
    output_declaration1247 output_declaration_instance1247();
    output_declaration1248 output_declaration_instance1248();
    output_declaration1249 output_declaration_instance1249();
    output_declaration1250 output_declaration_instance1250();
    output_declaration1251 output_declaration_instance1251();
    output_declaration1252 output_declaration_instance1252();
    output_declaration1253 output_declaration_instance1253();
    output_declaration1254 output_declaration_instance1254();
    output_declaration1255 output_declaration_instance1255();
    output_declaration1256 output_declaration_instance1256();
    output_declaration1257 output_declaration_instance1257();
    output_declaration1258 output_declaration_instance1258();
    output_declaration1259 output_declaration_instance1259();
    output_declaration1260 output_declaration_instance1260();
    output_declaration1261 output_declaration_instance1261();
    output_declaration1262 output_declaration_instance1262();
    output_declaration1263 output_declaration_instance1263();
    output_declaration1264 output_declaration_instance1264();
    output_declaration1265 output_declaration_instance1265();
    output_declaration1266 output_declaration_instance1266();
    output_declaration1267 output_declaration_instance1267();
    output_declaration1268 output_declaration_instance1268();
    output_declaration1269 output_declaration_instance1269();
    output_declaration1270 output_declaration_instance1270();
    output_declaration1271 output_declaration_instance1271();
    output_declaration1272 output_declaration_instance1272();
    output_declaration1273 output_declaration_instance1273();
    output_declaration1274 output_declaration_instance1274();
    output_declaration1275 output_declaration_instance1275();
    output_declaration1276 output_declaration_instance1276();
    output_declaration1277 output_declaration_instance1277();
    output_declaration1278 output_declaration_instance1278();
    output_declaration1279 output_declaration_instance1279();
    output_declaration1280 output_declaration_instance1280();
    output_declaration1281 output_declaration_instance1281();
    output_declaration1282 output_declaration_instance1282();
    output_declaration1283 output_declaration_instance1283();
    output_declaration1284 output_declaration_instance1284();
    output_declaration1285 output_declaration_instance1285();
    output_declaration1286 output_declaration_instance1286();
    output_declaration1287 output_declaration_instance1287();
    output_declaration1288 output_declaration_instance1288();
    output_declaration1289 output_declaration_instance1289();
    output_declaration1290 output_declaration_instance1290();
    output_declaration1291 output_declaration_instance1291();
    output_declaration1292 output_declaration_instance1292();
    output_declaration1293 output_declaration_instance1293();
    output_declaration1294 output_declaration_instance1294();
    output_declaration1295 output_declaration_instance1295();
    output_declaration1296 output_declaration_instance1296();
    output_declaration1297 output_declaration_instance1297();
    output_declaration1298 output_declaration_instance1298();
    output_declaration1299 output_declaration_instance1299();
    output_declaration1300 output_declaration_instance1300();
    output_declaration1301 output_declaration_instance1301();
    output_declaration1302 output_declaration_instance1302();
    output_declaration1303 output_declaration_instance1303();
    output_declaration1304 output_declaration_instance1304();
    output_declaration1305 output_declaration_instance1305();
    output_declaration1306 output_declaration_instance1306();
    output_declaration1307 output_declaration_instance1307();
    output_declaration1308 output_declaration_instance1308();
    output_declaration1309 output_declaration_instance1309();
    output_declaration1310 output_declaration_instance1310();
    output_declaration1311 output_declaration_instance1311();
    output_declaration1312 output_declaration_instance1312();
    output_declaration1313 output_declaration_instance1313();
    output_declaration1314 output_declaration_instance1314();
    output_declaration1315 output_declaration_instance1315();
    output_declaration1316 output_declaration_instance1316();
    output_declaration1317 output_declaration_instance1317();
    output_declaration1318 output_declaration_instance1318();
    output_declaration1319 output_declaration_instance1319();
    output_declaration1320 output_declaration_instance1320();
    output_declaration1321 output_declaration_instance1321();
    output_declaration1322 output_declaration_instance1322();
    output_declaration1323 output_declaration_instance1323();
    output_declaration1324 output_declaration_instance1324();
    output_declaration1325 output_declaration_instance1325();
    output_declaration1326 output_declaration_instance1326();
    output_declaration1327 output_declaration_instance1327();
    output_declaration1328 output_declaration_instance1328();
    output_declaration1329 output_declaration_instance1329();
    output_declaration1330 output_declaration_instance1330();
    output_declaration1331 output_declaration_instance1331();
    output_declaration1332 output_declaration_instance1332();
    output_declaration1333 output_declaration_instance1333();
    output_declaration1334 output_declaration_instance1334();
    output_declaration1335 output_declaration_instance1335();
    output_declaration1336 output_declaration_instance1336();
    output_declaration1337 output_declaration_instance1337();
    output_declaration1338 output_declaration_instance1338();
    output_declaration1339 output_declaration_instance1339();
    output_declaration1340 output_declaration_instance1340();
    output_declaration1341 output_declaration_instance1341();
    output_declaration1342 output_declaration_instance1342();
    output_declaration1343 output_declaration_instance1343();
    output_declaration1344 output_declaration_instance1344();
    output_declaration1345 output_declaration_instance1345();
    output_declaration1346 output_declaration_instance1346();
    output_declaration1347 output_declaration_instance1347();
    output_declaration1348 output_declaration_instance1348();
    output_declaration1349 output_declaration_instance1349();
    output_declaration1350 output_declaration_instance1350();
    output_declaration1351 output_declaration_instance1351();
    output_declaration1352 output_declaration_instance1352();
    output_declaration1353 output_declaration_instance1353();
    output_declaration1354 output_declaration_instance1354();
    output_declaration1355 output_declaration_instance1355();
    output_declaration1356 output_declaration_instance1356();
    output_declaration1357 output_declaration_instance1357();
    output_declaration1358 output_declaration_instance1358();
    output_declaration1359 output_declaration_instance1359();
    output_declaration1360 output_declaration_instance1360();
    output_declaration1361 output_declaration_instance1361();
    output_declaration1362 output_declaration_instance1362();
    output_declaration1363 output_declaration_instance1363();
    output_declaration1364 output_declaration_instance1364();
    output_declaration1365 output_declaration_instance1365();
    output_declaration1366 output_declaration_instance1366();
    output_declaration1367 output_declaration_instance1367();
    output_declaration1368 output_declaration_instance1368();
    output_declaration1369 output_declaration_instance1369();
    output_declaration1370 output_declaration_instance1370();
    output_declaration1371 output_declaration_instance1371();
    output_declaration1372 output_declaration_instance1372();
    output_declaration1373 output_declaration_instance1373();
    output_declaration1374 output_declaration_instance1374();
    output_declaration1375 output_declaration_instance1375();
    output_declaration1376 output_declaration_instance1376();
    output_declaration1377 output_declaration_instance1377();
    output_declaration1378 output_declaration_instance1378();
    output_declaration1379 output_declaration_instance1379();
    output_declaration1380 output_declaration_instance1380();
    output_declaration1381 output_declaration_instance1381();
    output_declaration1382 output_declaration_instance1382();
    output_declaration1383 output_declaration_instance1383();
    output_declaration1384 output_declaration_instance1384();
    output_declaration1385 output_declaration_instance1385();
    output_declaration1386 output_declaration_instance1386();
    output_declaration1387 output_declaration_instance1387();
    output_declaration1388 output_declaration_instance1388();
    output_declaration1389 output_declaration_instance1389();
    output_declaration1390 output_declaration_instance1390();
    output_declaration1391 output_declaration_instance1391();
    output_declaration1392 output_declaration_instance1392();
    output_declaration1393 output_declaration_instance1393();
    output_declaration1394 output_declaration_instance1394();
    output_declaration1395 output_declaration_instance1395();
    output_declaration1396 output_declaration_instance1396();
    output_declaration1397 output_declaration_instance1397();
    output_declaration1398 output_declaration_instance1398();
    output_declaration1399 output_declaration_instance1399();
    output_declaration1400 output_declaration_instance1400();
    output_declaration1401 output_declaration_instance1401();
    output_declaration1402 output_declaration_instance1402();
    output_declaration1403 output_declaration_instance1403();
    output_declaration1404 output_declaration_instance1404();
    output_declaration1405 output_declaration_instance1405();
    output_declaration1406 output_declaration_instance1406();
    output_declaration1407 output_declaration_instance1407();
    output_declaration1408 output_declaration_instance1408();
    output_declaration1409 output_declaration_instance1409();
    output_declaration1410 output_declaration_instance1410();
    output_declaration1411 output_declaration_instance1411();
    output_declaration1412 output_declaration_instance1412();
    output_declaration1413 output_declaration_instance1413();
    output_declaration1414 output_declaration_instance1414();
    output_declaration1415 output_declaration_instance1415();
    output_declaration1416 output_declaration_instance1416();
    output_declaration1417 output_declaration_instance1417();
    output_declaration1418 output_declaration_instance1418();
    output_declaration1419 output_declaration_instance1419();
    output_declaration1420 output_declaration_instance1420();
    output_declaration1421 output_declaration_instance1421();
    output_declaration1422 output_declaration_instance1422();
    output_declaration1423 output_declaration_instance1423();
    output_declaration1424 output_declaration_instance1424();
    output_declaration1425 output_declaration_instance1425();
    output_declaration1426 output_declaration_instance1426();
    output_declaration1427 output_declaration_instance1427();
    output_declaration1428 output_declaration_instance1428();
    output_declaration1429 output_declaration_instance1429();
    output_declaration1430 output_declaration_instance1430();
    output_declaration1431 output_declaration_instance1431();
    output_declaration1432 output_declaration_instance1432();
    output_declaration1433 output_declaration_instance1433();
    output_declaration1434 output_declaration_instance1434();
    output_declaration1435 output_declaration_instance1435();
    output_declaration1436 output_declaration_instance1436();
    output_declaration1437 output_declaration_instance1437();
    output_declaration1438 output_declaration_instance1438();
    output_declaration1439 output_declaration_instance1439();
    output_declaration1440 output_declaration_instance1440();
    output_declaration1441 output_declaration_instance1441();
    output_declaration1442 output_declaration_instance1442();
    output_declaration1443 output_declaration_instance1443();
    output_declaration1444 output_declaration_instance1444();
    output_declaration1445 output_declaration_instance1445();
    output_declaration1446 output_declaration_instance1446();
    output_declaration1447 output_declaration_instance1447();
    output_declaration1448 output_declaration_instance1448();
    output_declaration1449 output_declaration_instance1449();
    output_declaration1450 output_declaration_instance1450();
    output_declaration1451 output_declaration_instance1451();
    output_declaration1452 output_declaration_instance1452();
    output_declaration1453 output_declaration_instance1453();
    output_declaration1454 output_declaration_instance1454();
    output_declaration1455 output_declaration_instance1455();
    output_declaration1456 output_declaration_instance1456();
    output_declaration1457 output_declaration_instance1457();
    output_declaration1458 output_declaration_instance1458();
    output_declaration1459 output_declaration_instance1459();
    output_declaration1460 output_declaration_instance1460();
    output_declaration1461 output_declaration_instance1461();
    output_declaration1462 output_declaration_instance1462();
    output_declaration1463 output_declaration_instance1463();
    output_declaration1464 output_declaration_instance1464();
    output_declaration1465 output_declaration_instance1465();
    output_declaration1466 output_declaration_instance1466();
    output_declaration1467 output_declaration_instance1467();
    output_declaration1468 output_declaration_instance1468();
    output_declaration1469 output_declaration_instance1469();
    output_declaration1470 output_declaration_instance1470();
    output_declaration1471 output_declaration_instance1471();
    output_declaration1472 output_declaration_instance1472();
    output_declaration1473 output_declaration_instance1473();
    output_declaration1474 output_declaration_instance1474();
    output_declaration1475 output_declaration_instance1475();
    output_declaration1476 output_declaration_instance1476();
    output_declaration1477 output_declaration_instance1477();
    output_declaration1478 output_declaration_instance1478();
    output_declaration1479 output_declaration_instance1479();
    output_declaration1480 output_declaration_instance1480();
    output_declaration1481 output_declaration_instance1481();
    output_declaration1482 output_declaration_instance1482();
    output_declaration1483 output_declaration_instance1483();
    output_declaration1484 output_declaration_instance1484();
    output_declaration1485 output_declaration_instance1485();
    output_declaration1486 output_declaration_instance1486();
    output_declaration1487 output_declaration_instance1487();
    output_declaration1488 output_declaration_instance1488();
    output_declaration1489 output_declaration_instance1489();
    output_declaration1490 output_declaration_instance1490();
    output_declaration1491 output_declaration_instance1491();
    output_declaration1492 output_declaration_instance1492();
    output_declaration1493 output_declaration_instance1493();
    output_declaration1494 output_declaration_instance1494();
    output_declaration1495 output_declaration_instance1495();
    output_declaration1496 output_declaration_instance1496();
    output_declaration1497 output_declaration_instance1497();
    output_declaration1498 output_declaration_instance1498();
    output_declaration1499 output_declaration_instance1499();
    output_declaration1500 output_declaration_instance1500();
    output_declaration1501 output_declaration_instance1501();
    output_declaration1502 output_declaration_instance1502();
    output_declaration1503 output_declaration_instance1503();
    output_declaration1504 output_declaration_instance1504();
    output_declaration1505 output_declaration_instance1505();
    output_declaration1506 output_declaration_instance1506();
    output_declaration1507 output_declaration_instance1507();
    output_declaration1508 output_declaration_instance1508();
    output_declaration1509 output_declaration_instance1509();
    output_declaration1510 output_declaration_instance1510();
    output_declaration1511 output_declaration_instance1511();
    output_declaration1512 output_declaration_instance1512();
    output_declaration1513 output_declaration_instance1513();
    output_declaration1514 output_declaration_instance1514();
    output_declaration1515 output_declaration_instance1515();
    output_declaration1516 output_declaration_instance1516();
    output_declaration1517 output_declaration_instance1517();
    output_declaration1518 output_declaration_instance1518();
    output_declaration1519 output_declaration_instance1519();
    output_declaration1520 output_declaration_instance1520();
    output_declaration1521 output_declaration_instance1521();
    output_declaration1522 output_declaration_instance1522();
    output_declaration1523 output_declaration_instance1523();
    output_declaration1524 output_declaration_instance1524();
    output_declaration1525 output_declaration_instance1525();
    output_declaration1526 output_declaration_instance1526();
    output_declaration1527 output_declaration_instance1527();
    output_declaration1528 output_declaration_instance1528();
    output_declaration1529 output_declaration_instance1529();
    output_declaration1530 output_declaration_instance1530();
    output_declaration1531 output_declaration_instance1531();
    output_declaration1532 output_declaration_instance1532();
    output_declaration1533 output_declaration_instance1533();
    output_declaration1534 output_declaration_instance1534();
    output_declaration1535 output_declaration_instance1535();
    output_declaration1536 output_declaration_instance1536();
    output_declaration1537 output_declaration_instance1537();
    output_declaration1538 output_declaration_instance1538();
    output_declaration1539 output_declaration_instance1539();
    output_declaration1540 output_declaration_instance1540();
    output_declaration1541 output_declaration_instance1541();
    output_declaration1542 output_declaration_instance1542();
    output_declaration1543 output_declaration_instance1543();
    output_declaration1544 output_declaration_instance1544();
    output_declaration1545 output_declaration_instance1545();
    output_declaration1546 output_declaration_instance1546();
    output_declaration1547 output_declaration_instance1547();
    output_declaration1548 output_declaration_instance1548();
    output_declaration1549 output_declaration_instance1549();
    output_declaration1550 output_declaration_instance1550();
    output_declaration1551 output_declaration_instance1551();
    output_declaration1552 output_declaration_instance1552();
    output_declaration1553 output_declaration_instance1553();
    output_declaration1554 output_declaration_instance1554();
    output_declaration1555 output_declaration_instance1555();
    output_declaration1556 output_declaration_instance1556();
    output_declaration1557 output_declaration_instance1557();
    output_declaration1558 output_declaration_instance1558();
    output_declaration1559 output_declaration_instance1559();
    output_declaration1560 output_declaration_instance1560();
    output_declaration1561 output_declaration_instance1561();
    output_declaration1562 output_declaration_instance1562();
    output_declaration1563 output_declaration_instance1563();
    output_declaration1564 output_declaration_instance1564();
    output_declaration1565 output_declaration_instance1565();
    output_declaration1566 output_declaration_instance1566();
    output_declaration1567 output_declaration_instance1567();
    output_declaration1568 output_declaration_instance1568();
    output_declaration1569 output_declaration_instance1569();
    output_declaration1570 output_declaration_instance1570();
    output_declaration1571 output_declaration_instance1571();
    output_declaration1572 output_declaration_instance1572();
    output_declaration1573 output_declaration_instance1573();
    output_declaration1574 output_declaration_instance1574();
    output_declaration1575 output_declaration_instance1575();
    output_declaration1576 output_declaration_instance1576();
    output_declaration1577 output_declaration_instance1577();
    output_declaration1578 output_declaration_instance1578();
    output_declaration1579 output_declaration_instance1579();
    output_declaration1580 output_declaration_instance1580();
    output_declaration1581 output_declaration_instance1581();
    output_declaration1582 output_declaration_instance1582();
    output_declaration1583 output_declaration_instance1583();
    output_declaration1584 output_declaration_instance1584();
    output_declaration1585 output_declaration_instance1585();
    output_declaration1586 output_declaration_instance1586();
    output_declaration1587 output_declaration_instance1587();
    output_declaration1588 output_declaration_instance1588();
    output_declaration1589 output_declaration_instance1589();
    output_declaration1590 output_declaration_instance1590();
    output_declaration1591 output_declaration_instance1591();
    output_declaration1592 output_declaration_instance1592();
    output_declaration1593 output_declaration_instance1593();
    output_declaration1594 output_declaration_instance1594();
    output_declaration1595 output_declaration_instance1595();
    output_declaration1596 output_declaration_instance1596();
    output_declaration1597 output_declaration_instance1597();
    output_declaration1598 output_declaration_instance1598();
    output_declaration1599 output_declaration_instance1599();
    output_declaration1600 output_declaration_instance1600();
    output_declaration1601 output_declaration_instance1601();
    output_declaration1602 output_declaration_instance1602();
    output_declaration1603 output_declaration_instance1603();
    output_declaration1604 output_declaration_instance1604();
    output_declaration1605 output_declaration_instance1605();
    output_declaration1606 output_declaration_instance1606();
    output_declaration1607 output_declaration_instance1607();
    output_declaration1608 output_declaration_instance1608();
    output_declaration1609 output_declaration_instance1609();
    output_declaration1610 output_declaration_instance1610();
    output_declaration1611 output_declaration_instance1611();
    output_declaration1612 output_declaration_instance1612();
    output_declaration1613 output_declaration_instance1613();
    output_declaration1614 output_declaration_instance1614();
    output_declaration1615 output_declaration_instance1615();
    output_declaration1616 output_declaration_instance1616();
    output_declaration1617 output_declaration_instance1617();
    output_declaration1618 output_declaration_instance1618();
    output_declaration1619 output_declaration_instance1619();
    output_declaration1620 output_declaration_instance1620();
    output_declaration1621 output_declaration_instance1621();
    output_declaration1622 output_declaration_instance1622();
    output_declaration1623 output_declaration_instance1623();
    output_declaration1624 output_declaration_instance1624();
    output_declaration1625 output_declaration_instance1625();
    output_declaration1626 output_declaration_instance1626();
    output_declaration1627 output_declaration_instance1627();
    output_declaration1628 output_declaration_instance1628();
    output_declaration1629 output_declaration_instance1629();
    output_declaration1630 output_declaration_instance1630();
    output_declaration1631 output_declaration_instance1631();
    output_declaration1632 output_declaration_instance1632();
    output_declaration1633 output_declaration_instance1633();
    output_declaration1634 output_declaration_instance1634();
    output_declaration1635 output_declaration_instance1635();
    output_declaration1636 output_declaration_instance1636();
    output_declaration1637 output_declaration_instance1637();
    output_declaration1638 output_declaration_instance1638();
    output_declaration1639 output_declaration_instance1639();
    output_declaration1640 output_declaration_instance1640();
    output_declaration1641 output_declaration_instance1641();
    output_declaration1642 output_declaration_instance1642();
    output_declaration1643 output_declaration_instance1643();
    output_declaration1644 output_declaration_instance1644();
    output_declaration1645 output_declaration_instance1645();
    output_declaration1646 output_declaration_instance1646();
    output_declaration1647 output_declaration_instance1647();
    output_declaration1648 output_declaration_instance1648();
    output_declaration1649 output_declaration_instance1649();
    output_declaration1650 output_declaration_instance1650();
    output_declaration1651 output_declaration_instance1651();
    output_declaration1652 output_declaration_instance1652();
    output_declaration1653 output_declaration_instance1653();
    output_declaration1654 output_declaration_instance1654();
    output_declaration1655 output_declaration_instance1655();
    output_declaration1656 output_declaration_instance1656();
    output_declaration1657 output_declaration_instance1657();
    output_declaration1658 output_declaration_instance1658();
    output_declaration1659 output_declaration_instance1659();
    output_declaration1660 output_declaration_instance1660();
    output_declaration1661 output_declaration_instance1661();
    output_declaration1662 output_declaration_instance1662();
    output_declaration1663 output_declaration_instance1663();
    output_declaration1664 output_declaration_instance1664();
    output_declaration1665 output_declaration_instance1665();
    output_declaration1666 output_declaration_instance1666();
    output_declaration1667 output_declaration_instance1667();
    output_declaration1668 output_declaration_instance1668();
    output_declaration1669 output_declaration_instance1669();
    output_declaration1670 output_declaration_instance1670();
    output_declaration1671 output_declaration_instance1671();
    output_declaration1672 output_declaration_instance1672();
    output_declaration1673 output_declaration_instance1673();
    output_declaration1674 output_declaration_instance1674();
    output_declaration1675 output_declaration_instance1675();
    output_declaration1676 output_declaration_instance1676();
    output_declaration1677 output_declaration_instance1677();
    output_declaration1678 output_declaration_instance1678();
    output_declaration1679 output_declaration_instance1679();
    output_declaration1680 output_declaration_instance1680();
    output_declaration1681 output_declaration_instance1681();
    output_declaration1682 output_declaration_instance1682();
    output_declaration1683 output_declaration_instance1683();
    output_declaration1684 output_declaration_instance1684();
    output_declaration1685 output_declaration_instance1685();
    output_declaration1686 output_declaration_instance1686();
    output_declaration1687 output_declaration_instance1687();
    output_declaration1688 output_declaration_instance1688();
    output_declaration1689 output_declaration_instance1689();
    output_declaration1690 output_declaration_instance1690();
    output_declaration1691 output_declaration_instance1691();
    output_declaration1692 output_declaration_instance1692();
    output_declaration1693 output_declaration_instance1693();
    output_declaration1694 output_declaration_instance1694();
    output_declaration1695 output_declaration_instance1695();
    output_declaration1696 output_declaration_instance1696();
    output_declaration1697 output_declaration_instance1697();
    output_declaration1698 output_declaration_instance1698();
    output_declaration1699 output_declaration_instance1699();
    output_declaration1700 output_declaration_instance1700();
    output_declaration1701 output_declaration_instance1701();
    output_declaration1702 output_declaration_instance1702();
    output_declaration1703 output_declaration_instance1703();
    output_declaration1704 output_declaration_instance1704();
    output_declaration1705 output_declaration_instance1705();
    output_declaration1706 output_declaration_instance1706();
    output_declaration1707 output_declaration_instance1707();
    output_declaration1708 output_declaration_instance1708();
    output_declaration1709 output_declaration_instance1709();
    output_declaration1710 output_declaration_instance1710();
    output_declaration1711 output_declaration_instance1711();
    output_declaration1712 output_declaration_instance1712();
    output_declaration1713 output_declaration_instance1713();
    output_declaration1714 output_declaration_instance1714();
    output_declaration1715 output_declaration_instance1715();
    output_declaration1716 output_declaration_instance1716();
    output_declaration1717 output_declaration_instance1717();
    output_declaration1718 output_declaration_instance1718();
    output_declaration1719 output_declaration_instance1719();
    output_declaration1720 output_declaration_instance1720();
    output_declaration1721 output_declaration_instance1721();
    output_declaration1722 output_declaration_instance1722();
    output_declaration1723 output_declaration_instance1723();
    output_declaration1724 output_declaration_instance1724();
    output_declaration1725 output_declaration_instance1725();
    output_declaration1726 output_declaration_instance1726();
    output_declaration1727 output_declaration_instance1727();
    output_declaration1728 output_declaration_instance1728();
    output_declaration1729 output_declaration_instance1729();
    output_declaration1730 output_declaration_instance1730();
    output_declaration1731 output_declaration_instance1731();
    output_declaration1732 output_declaration_instance1732();
    output_declaration1733 output_declaration_instance1733();
    output_declaration1734 output_declaration_instance1734();
    output_declaration1735 output_declaration_instance1735();
    output_declaration1736 output_declaration_instance1736();
    output_declaration1737 output_declaration_instance1737();
    output_declaration1738 output_declaration_instance1738();
    output_declaration1739 output_declaration_instance1739();
    output_declaration1740 output_declaration_instance1740();
    output_declaration1741 output_declaration_instance1741();
    output_declaration1742 output_declaration_instance1742();
    output_declaration1743 output_declaration_instance1743();
    output_declaration1744 output_declaration_instance1744();
    output_declaration1745 output_declaration_instance1745();
    output_declaration1746 output_declaration_instance1746();
    output_declaration1747 output_declaration_instance1747();
    output_declaration1748 output_declaration_instance1748();
    output_declaration1749 output_declaration_instance1749();
    output_declaration1750 output_declaration_instance1750();
    output_declaration1751 output_declaration_instance1751();
    output_declaration1752 output_declaration_instance1752();
    output_declaration1753 output_declaration_instance1753();
    output_declaration1754 output_declaration_instance1754();
    output_declaration1755 output_declaration_instance1755();
    output_declaration1756 output_declaration_instance1756();
    output_declaration1757 output_declaration_instance1757();
    output_declaration1758 output_declaration_instance1758();
    output_declaration1759 output_declaration_instance1759();
    output_declaration1760 output_declaration_instance1760();
    output_declaration1761 output_declaration_instance1761();
    output_declaration1762 output_declaration_instance1762();
    output_declaration1763 output_declaration_instance1763();
    output_declaration1764 output_declaration_instance1764();
    output_declaration1765 output_declaration_instance1765();
    output_declaration1766 output_declaration_instance1766();
    output_declaration1767 output_declaration_instance1767();
    output_declaration1768 output_declaration_instance1768();
    output_declaration1769 output_declaration_instance1769();
    output_declaration1770 output_declaration_instance1770();
    output_declaration1771 output_declaration_instance1771();
    output_declaration1772 output_declaration_instance1772();
    output_declaration1773 output_declaration_instance1773();
    output_declaration1774 output_declaration_instance1774();
    output_declaration1775 output_declaration_instance1775();
    output_declaration1776 output_declaration_instance1776();
    output_declaration1777 output_declaration_instance1777();
    output_declaration1778 output_declaration_instance1778();
    output_declaration1779 output_declaration_instance1779();
    output_declaration1780 output_declaration_instance1780();
    output_declaration1781 output_declaration_instance1781();
    output_declaration1782 output_declaration_instance1782();
    output_declaration1783 output_declaration_instance1783();
    output_declaration1784 output_declaration_instance1784();
    output_declaration1785 output_declaration_instance1785();
    output_declaration1786 output_declaration_instance1786();
    output_declaration1787 output_declaration_instance1787();
    output_declaration1788 output_declaration_instance1788();
    output_declaration1789 output_declaration_instance1789();
    output_declaration1790 output_declaration_instance1790();
    output_declaration1791 output_declaration_instance1791();
    output_declaration1792 output_declaration_instance1792();
    output_declaration1793 output_declaration_instance1793();
    output_declaration1794 output_declaration_instance1794();
    output_declaration1795 output_declaration_instance1795();
    output_declaration1796 output_declaration_instance1796();
    output_declaration1797 output_declaration_instance1797();
    output_declaration1798 output_declaration_instance1798();
    output_declaration1799 output_declaration_instance1799();
    output_declaration1800 output_declaration_instance1800();
    output_declaration1801 output_declaration_instance1801();
    output_declaration1802 output_declaration_instance1802();
    output_declaration1803 output_declaration_instance1803();
    output_declaration1804 output_declaration_instance1804();
    output_declaration1805 output_declaration_instance1805();
    output_declaration1806 output_declaration_instance1806();
    output_declaration1807 output_declaration_instance1807();
    output_declaration1808 output_declaration_instance1808();
    output_declaration1809 output_declaration_instance1809();
    output_declaration1810 output_declaration_instance1810();
    output_declaration1811 output_declaration_instance1811();
    output_declaration1812 output_declaration_instance1812();
    output_declaration1813 output_declaration_instance1813();
    output_declaration1814 output_declaration_instance1814();
    output_declaration1815 output_declaration_instance1815();
    output_declaration1816 output_declaration_instance1816();
    output_declaration1817 output_declaration_instance1817();
    output_declaration1818 output_declaration_instance1818();
    output_declaration1819 output_declaration_instance1819();
    output_declaration1820 output_declaration_instance1820();
    output_declaration1821 output_declaration_instance1821();
    output_declaration1822 output_declaration_instance1822();
    output_declaration1823 output_declaration_instance1823();
    output_declaration1824 output_declaration_instance1824();
    output_declaration1825 output_declaration_instance1825();
    output_declaration1826 output_declaration_instance1826();
    output_declaration1827 output_declaration_instance1827();
    output_declaration1828 output_declaration_instance1828();
    output_declaration1829 output_declaration_instance1829();
    output_declaration1830 output_declaration_instance1830();
    output_declaration1831 output_declaration_instance1831();
    output_declaration1832 output_declaration_instance1832();
    output_declaration1833 output_declaration_instance1833();
    output_declaration1834 output_declaration_instance1834();
    output_declaration1835 output_declaration_instance1835();
    output_declaration1836 output_declaration_instance1836();
    output_declaration1837 output_declaration_instance1837();
    output_declaration1838 output_declaration_instance1838();
    output_declaration1839 output_declaration_instance1839();
    output_declaration1840 output_declaration_instance1840();
    output_declaration1841 output_declaration_instance1841();
    output_declaration1842 output_declaration_instance1842();
    output_declaration1843 output_declaration_instance1843();
    output_declaration1844 output_declaration_instance1844();
    output_declaration1845 output_declaration_instance1845();
    output_declaration1846 output_declaration_instance1846();
    output_declaration1847 output_declaration_instance1847();
    output_declaration1848 output_declaration_instance1848();
    output_declaration1849 output_declaration_instance1849();
    output_declaration1850 output_declaration_instance1850();
    output_declaration1851 output_declaration_instance1851();
    output_declaration1852 output_declaration_instance1852();
    output_declaration1853 output_declaration_instance1853();
    output_declaration1854 output_declaration_instance1854();
    output_declaration1855 output_declaration_instance1855();
    output_declaration1856 output_declaration_instance1856();
    output_declaration1857 output_declaration_instance1857();
    output_declaration1858 output_declaration_instance1858();
    output_declaration1859 output_declaration_instance1859();
    output_declaration1860 output_declaration_instance1860();
    output_declaration1861 output_declaration_instance1861();
    output_declaration1862 output_declaration_instance1862();
    output_declaration1863 output_declaration_instance1863();
    output_declaration1864 output_declaration_instance1864();
    output_declaration1865 output_declaration_instance1865();
    output_declaration1866 output_declaration_instance1866();
    output_declaration1867 output_declaration_instance1867();
    output_declaration1868 output_declaration_instance1868();
    output_declaration1869 output_declaration_instance1869();
    output_declaration1870 output_declaration_instance1870();
    output_declaration1871 output_declaration_instance1871();
    output_declaration1872 output_declaration_instance1872();
    output_declaration1873 output_declaration_instance1873();
    output_declaration1874 output_declaration_instance1874();
    output_declaration1875 output_declaration_instance1875();
    output_declaration1876 output_declaration_instance1876();
    output_declaration1877 output_declaration_instance1877();
    output_declaration1878 output_declaration_instance1878();
    output_declaration1879 output_declaration_instance1879();
    output_declaration1880 output_declaration_instance1880();
    output_declaration1881 output_declaration_instance1881();
    output_declaration1882 output_declaration_instance1882();
    output_declaration1883 output_declaration_instance1883();
    output_declaration1884 output_declaration_instance1884();
    output_declaration1885 output_declaration_instance1885();
    output_declaration1886 output_declaration_instance1886();
    output_declaration1887 output_declaration_instance1887();
    output_declaration1888 output_declaration_instance1888();
    output_declaration1889 output_declaration_instance1889();
    output_declaration1890 output_declaration_instance1890();
    output_declaration1891 output_declaration_instance1891();
    output_declaration1892 output_declaration_instance1892();
    output_declaration1893 output_declaration_instance1893();
    output_declaration1894 output_declaration_instance1894();
    output_declaration1895 output_declaration_instance1895();
    output_declaration1896 output_declaration_instance1896();
    output_declaration1897 output_declaration_instance1897();
    output_declaration1898 output_declaration_instance1898();
    output_declaration1899 output_declaration_instance1899();
    output_declaration1900 output_declaration_instance1900();
    output_declaration1901 output_declaration_instance1901();
    output_declaration1902 output_declaration_instance1902();
    output_declaration1903 output_declaration_instance1903();
    output_declaration1904 output_declaration_instance1904();
    output_declaration1905 output_declaration_instance1905();
    output_declaration1906 output_declaration_instance1906();
    output_declaration1907 output_declaration_instance1907();
    output_declaration1908 output_declaration_instance1908();
    output_declaration1909 output_declaration_instance1909();
    output_declaration1910 output_declaration_instance1910();
    output_declaration1911 output_declaration_instance1911();
    output_declaration1912 output_declaration_instance1912();
    output_declaration1913 output_declaration_instance1913();
    output_declaration1914 output_declaration_instance1914();
    output_declaration1915 output_declaration_instance1915();
    output_declaration1916 output_declaration_instance1916();
    output_declaration1917 output_declaration_instance1917();
    output_declaration1918 output_declaration_instance1918();
    output_declaration1919 output_declaration_instance1919();
    output_declaration1920 output_declaration_instance1920();
    output_declaration1921 output_declaration_instance1921();
    output_declaration1922 output_declaration_instance1922();
    output_declaration1923 output_declaration_instance1923();
    output_declaration1924 output_declaration_instance1924();
    output_declaration1925 output_declaration_instance1925();
    output_declaration1926 output_declaration_instance1926();
    output_declaration1927 output_declaration_instance1927();
    output_declaration1928 output_declaration_instance1928();
    output_declaration1929 output_declaration_instance1929();
    output_declaration1930 output_declaration_instance1930();
    output_declaration1931 output_declaration_instance1931();
    output_declaration1932 output_declaration_instance1932();
    output_declaration1933 output_declaration_instance1933();
    output_declaration1934 output_declaration_instance1934();
    output_declaration1935 output_declaration_instance1935();
    output_declaration1936 output_declaration_instance1936();
    output_declaration1937 output_declaration_instance1937();
    output_declaration1938 output_declaration_instance1938();
    output_declaration1939 output_declaration_instance1939();
    output_declaration1940 output_declaration_instance1940();
    output_declaration1941 output_declaration_instance1941();
    output_declaration1942 output_declaration_instance1942();
    output_declaration1943 output_declaration_instance1943();
    output_declaration1944 output_declaration_instance1944();
    output_declaration1945 output_declaration_instance1945();
    output_declaration1946 output_declaration_instance1946();
    output_declaration1947 output_declaration_instance1947();
    output_declaration1948 output_declaration_instance1948();
    output_declaration1949 output_declaration_instance1949();
    output_declaration1950 output_declaration_instance1950();
    output_declaration1951 output_declaration_instance1951();
    output_declaration1952 output_declaration_instance1952();
    output_declaration1953 output_declaration_instance1953();
    output_declaration1954 output_declaration_instance1954();
    output_declaration1955 output_declaration_instance1955();
    output_declaration1956 output_declaration_instance1956();
    output_declaration1957 output_declaration_instance1957();
    output_declaration1958 output_declaration_instance1958();
    output_declaration1959 output_declaration_instance1959();
    output_declaration1960 output_declaration_instance1960();
    output_declaration1961 output_declaration_instance1961();
    output_declaration1962 output_declaration_instance1962();
    output_declaration1963 output_declaration_instance1963();
    output_declaration1964 output_declaration_instance1964();
    output_declaration1965 output_declaration_instance1965();
    output_declaration1966 output_declaration_instance1966();
    output_declaration1967 output_declaration_instance1967();
    output_declaration1968 output_declaration_instance1968();
    output_declaration1969 output_declaration_instance1969();
    output_declaration1970 output_declaration_instance1970();
    output_declaration1971 output_declaration_instance1971();
    output_declaration1972 output_declaration_instance1972();
    output_declaration1973 output_declaration_instance1973();
    output_declaration1974 output_declaration_instance1974();
    output_declaration1975 output_declaration_instance1975();
    output_declaration1976 output_declaration_instance1976();
    output_declaration1977 output_declaration_instance1977();
    output_declaration1978 output_declaration_instance1978();
    output_declaration1979 output_declaration_instance1979();
    output_declaration1980 output_declaration_instance1980();
    output_declaration1981 output_declaration_instance1981();
    output_declaration1982 output_declaration_instance1982();
    output_declaration1983 output_declaration_instance1983();
    output_declaration1984 output_declaration_instance1984();
    output_declaration1985 output_declaration_instance1985();
    output_declaration1986 output_declaration_instance1986();
    output_declaration1987 output_declaration_instance1987();
    output_declaration1988 output_declaration_instance1988();
    output_declaration1989 output_declaration_instance1989();
    output_declaration1990 output_declaration_instance1990();
    output_declaration1991 output_declaration_instance1991();
    output_declaration1992 output_declaration_instance1992();
    output_declaration1993 output_declaration_instance1993();
    output_declaration1994 output_declaration_instance1994();
    output_declaration1995 output_declaration_instance1995();
    output_declaration1996 output_declaration_instance1996();
    output_declaration1997 output_declaration_instance1997();
    output_declaration1998 output_declaration_instance1998();
    output_declaration1999 output_declaration_instance1999();
    output_declaration2000 output_declaration_instance2000();
    output_declaration2001 output_declaration_instance2001();
    output_declaration2002 output_declaration_instance2002();
    output_declaration2003 output_declaration_instance2003();
    output_declaration2004 output_declaration_instance2004();
    output_declaration2005 output_declaration_instance2005();
    output_declaration2006 output_declaration_instance2006();
    output_declaration2007 output_declaration_instance2007();
    output_declaration2008 output_declaration_instance2008();
    output_declaration2009 output_declaration_instance2009();
    output_declaration2010 output_declaration_instance2010();
    output_declaration2011 output_declaration_instance2011();
    output_declaration2012 output_declaration_instance2012();
    output_declaration2013 output_declaration_instance2013();
    output_declaration2014 output_declaration_instance2014();
    output_declaration2015 output_declaration_instance2015();
    output_declaration2016 output_declaration_instance2016();
    output_declaration2017 output_declaration_instance2017();
    output_declaration2018 output_declaration_instance2018();
    output_declaration2019 output_declaration_instance2019();
    output_declaration2020 output_declaration_instance2020();
    output_declaration2021 output_declaration_instance2021();
    output_declaration2022 output_declaration_instance2022();
    output_declaration2023 output_declaration_instance2023();
    output_declaration2024 output_declaration_instance2024();
    output_declaration2025 output_declaration_instance2025();
    output_declaration2026 output_declaration_instance2026();
    output_declaration2027 output_declaration_instance2027();
    output_declaration2028 output_declaration_instance2028();
    output_declaration2029 output_declaration_instance2029();
    output_declaration2030 output_declaration_instance2030();
    output_declaration2031 output_declaration_instance2031();
    output_declaration2032 output_declaration_instance2032();
    output_declaration2033 output_declaration_instance2033();
    output_declaration2034 output_declaration_instance2034();
    output_declaration2035 output_declaration_instance2035();
    output_declaration2036 output_declaration_instance2036();
    output_declaration2037 output_declaration_instance2037();
    output_declaration2038 output_declaration_instance2038();
    output_declaration2039 output_declaration_instance2039();
    output_declaration2040 output_declaration_instance2040();
    output_declaration2041 output_declaration_instance2041();
    output_declaration2042 output_declaration_instance2042();
    output_declaration2043 output_declaration_instance2043();
    output_declaration2044 output_declaration_instance2044();
    output_declaration2045 output_declaration_instance2045();
    output_declaration2046 output_declaration_instance2046();
    output_declaration2047 output_declaration_instance2047();
    output_declaration2048 output_declaration_instance2048();
    output_declaration2049 output_declaration_instance2049();
    output_declaration2050 output_declaration_instance2050();
    output_declaration2051 output_declaration_instance2051();
    output_declaration2052 output_declaration_instance2052();
    output_declaration2053 output_declaration_instance2053();
    output_declaration2054 output_declaration_instance2054();
    output_declaration2055 output_declaration_instance2055();
    output_declaration2056 output_declaration_instance2056();
    output_declaration2057 output_declaration_instance2057();
    output_declaration2058 output_declaration_instance2058();
    output_declaration2059 output_declaration_instance2059();
    output_declaration2060 output_declaration_instance2060();
    output_declaration2061 output_declaration_instance2061();
    output_declaration2062 output_declaration_instance2062();
    output_declaration2063 output_declaration_instance2063();
    output_declaration2064 output_declaration_instance2064();
    output_declaration2065 output_declaration_instance2065();
    output_declaration2066 output_declaration_instance2066();
    output_declaration2067 output_declaration_instance2067();
    output_declaration2068 output_declaration_instance2068();
    output_declaration2069 output_declaration_instance2069();
    output_declaration2070 output_declaration_instance2070();
    output_declaration2071 output_declaration_instance2071();
    output_declaration2072 output_declaration_instance2072();
    output_declaration2073 output_declaration_instance2073();
    output_declaration2074 output_declaration_instance2074();
    output_declaration2075 output_declaration_instance2075();
    output_declaration2076 output_declaration_instance2076();
    output_declaration2077 output_declaration_instance2077();
    output_declaration2078 output_declaration_instance2078();
    output_declaration2079 output_declaration_instance2079();
    output_declaration2080 output_declaration_instance2080();
    output_declaration2081 output_declaration_instance2081();
    output_declaration2082 output_declaration_instance2082();
    output_declaration2083 output_declaration_instance2083();
    output_declaration2084 output_declaration_instance2084();
    output_declaration2085 output_declaration_instance2085();
    output_declaration2086 output_declaration_instance2086();
    output_declaration2087 output_declaration_instance2087();
    output_declaration2088 output_declaration_instance2088();
    output_declaration2089 output_declaration_instance2089();
    output_declaration2090 output_declaration_instance2090();
    output_declaration2091 output_declaration_instance2091();
    output_declaration2092 output_declaration_instance2092();
    output_declaration2093 output_declaration_instance2093();
    output_declaration2094 output_declaration_instance2094();
    output_declaration2095 output_declaration_instance2095();
    output_declaration2096 output_declaration_instance2096();
    output_declaration2097 output_declaration_instance2097();
    output_declaration2098 output_declaration_instance2098();
    output_declaration2099 output_declaration_instance2099();
    output_declaration2100 output_declaration_instance2100();
    output_declaration2101 output_declaration_instance2101();
    output_declaration2102 output_declaration_instance2102();
    output_declaration2103 output_declaration_instance2103();
    output_declaration2104 output_declaration_instance2104();
    output_declaration2105 output_declaration_instance2105();
    output_declaration2106 output_declaration_instance2106();
    output_declaration2107 output_declaration_instance2107();
    output_declaration2108 output_declaration_instance2108();
    output_declaration2109 output_declaration_instance2109();
    output_declaration2110 output_declaration_instance2110();
    output_declaration2111 output_declaration_instance2111();
    output_declaration2112 output_declaration_instance2112();
    output_declaration2113 output_declaration_instance2113();
    output_declaration2114 output_declaration_instance2114();
    output_declaration2115 output_declaration_instance2115();
    output_declaration2116 output_declaration_instance2116();
    output_declaration2117 output_declaration_instance2117();
    output_declaration2118 output_declaration_instance2118();
    output_declaration2119 output_declaration_instance2119();
    output_declaration2120 output_declaration_instance2120();
    output_declaration2121 output_declaration_instance2121();
    output_declaration2122 output_declaration_instance2122();
    output_declaration2123 output_declaration_instance2123();
    output_declaration2124 output_declaration_instance2124();
    output_declaration2125 output_declaration_instance2125();
    output_declaration2126 output_declaration_instance2126();
    output_declaration2127 output_declaration_instance2127();
    output_declaration2128 output_declaration_instance2128();
    output_declaration2129 output_declaration_instance2129();
    output_declaration2130 output_declaration_instance2130();
    output_declaration2131 output_declaration_instance2131();
    output_declaration2132 output_declaration_instance2132();
    output_declaration2133 output_declaration_instance2133();
    output_declaration2134 output_declaration_instance2134();
    output_declaration2135 output_declaration_instance2135();
    output_declaration2136 output_declaration_instance2136();
    output_declaration2137 output_declaration_instance2137();
    output_declaration2138 output_declaration_instance2138();
    output_declaration2139 output_declaration_instance2139();
    output_declaration2140 output_declaration_instance2140();
    output_declaration2141 output_declaration_instance2141();
    output_declaration2142 output_declaration_instance2142();
    output_declaration2143 output_declaration_instance2143();
    output_declaration2144 output_declaration_instance2144();
    output_declaration2145 output_declaration_instance2145();
    output_declaration2146 output_declaration_instance2146();
    output_declaration2147 output_declaration_instance2147();
    output_declaration2148 output_declaration_instance2148();
    output_declaration2149 output_declaration_instance2149();
    output_declaration2150 output_declaration_instance2150();
    output_declaration2151 output_declaration_instance2151();
    output_declaration2152 output_declaration_instance2152();
    output_declaration2153 output_declaration_instance2153();
    output_declaration2154 output_declaration_instance2154();
    output_declaration2155 output_declaration_instance2155();
    output_declaration2156 output_declaration_instance2156();
    output_declaration2157 output_declaration_instance2157();
    output_declaration2158 output_declaration_instance2158();
    output_declaration2159 output_declaration_instance2159();
    output_declaration2160 output_declaration_instance2160();
    output_declaration2161 output_declaration_instance2161();
    output_declaration2162 output_declaration_instance2162();
    output_declaration2163 output_declaration_instance2163();
    output_declaration2164 output_declaration_instance2164();
    output_declaration2165 output_declaration_instance2165();
    output_declaration2166 output_declaration_instance2166();
    output_declaration2167 output_declaration_instance2167();
    output_declaration2168 output_declaration_instance2168();
    output_declaration2169 output_declaration_instance2169();
    output_declaration2170 output_declaration_instance2170();
    output_declaration2171 output_declaration_instance2171();
    output_declaration2172 output_declaration_instance2172();
    output_declaration2173 output_declaration_instance2173();
    output_declaration2174 output_declaration_instance2174();
    output_declaration2175 output_declaration_instance2175();
    output_declaration2176 output_declaration_instance2176();
    output_declaration2177 output_declaration_instance2177();
    output_declaration2178 output_declaration_instance2178();
    output_declaration2179 output_declaration_instance2179();
    output_declaration2180 output_declaration_instance2180();
    output_declaration2181 output_declaration_instance2181();
    output_declaration2182 output_declaration_instance2182();
    output_declaration2183 output_declaration_instance2183();
    output_declaration2184 output_declaration_instance2184();
    output_declaration2185 output_declaration_instance2185();
    output_declaration2186 output_declaration_instance2186();
    output_declaration2187 output_declaration_instance2187();
    output_declaration2188 output_declaration_instance2188();
    output_declaration2189 output_declaration_instance2189();
    output_declaration2190 output_declaration_instance2190();
    output_declaration2191 output_declaration_instance2191();
    output_declaration2192 output_declaration_instance2192();
    output_declaration2193 output_declaration_instance2193();
    output_declaration2194 output_declaration_instance2194();
    output_declaration2195 output_declaration_instance2195();
    output_declaration2196 output_declaration_instance2196();
    output_declaration2197 output_declaration_instance2197();
    output_declaration2198 output_declaration_instance2198();
    output_declaration2199 output_declaration_instance2199();
    output_declaration2200 output_declaration_instance2200();
    output_declaration2201 output_declaration_instance2201();
    output_declaration2202 output_declaration_instance2202();
    output_declaration2203 output_declaration_instance2203();
    output_declaration2204 output_declaration_instance2204();
    output_declaration2205 output_declaration_instance2205();
    output_declaration2206 output_declaration_instance2206();
    output_declaration2207 output_declaration_instance2207();
    output_declaration2208 output_declaration_instance2208();
    output_declaration2209 output_declaration_instance2209();
    output_declaration2210 output_declaration_instance2210();
    output_declaration2211 output_declaration_instance2211();
    output_declaration2212 output_declaration_instance2212();
    output_declaration2213 output_declaration_instance2213();
    output_declaration2214 output_declaration_instance2214();
    output_declaration2215 output_declaration_instance2215();
    output_declaration2216 output_declaration_instance2216();
    output_declaration2217 output_declaration_instance2217();
    output_declaration2218 output_declaration_instance2218();
    output_declaration2219 output_declaration_instance2219();
    output_declaration2220 output_declaration_instance2220();
    output_declaration2221 output_declaration_instance2221();
    output_declaration2222 output_declaration_instance2222();
    output_declaration2223 output_declaration_instance2223();
    output_declaration2224 output_declaration_instance2224();
    output_declaration2225 output_declaration_instance2225();
    output_declaration2226 output_declaration_instance2226();
    output_declaration2227 output_declaration_instance2227();
    output_declaration2228 output_declaration_instance2228();
    output_declaration2229 output_declaration_instance2229();
    output_declaration2230 output_declaration_instance2230();
    output_declaration2231 output_declaration_instance2231();
    output_declaration2232 output_declaration_instance2232();
    output_declaration2233 output_declaration_instance2233();
    output_declaration2234 output_declaration_instance2234();
    output_declaration2235 output_declaration_instance2235();
    output_declaration2236 output_declaration_instance2236();
    output_declaration2237 output_declaration_instance2237();
    output_declaration2238 output_declaration_instance2238();
    output_declaration2239 output_declaration_instance2239();
    output_declaration2240 output_declaration_instance2240();
    output_declaration2241 output_declaration_instance2241();
    output_declaration2242 output_declaration_instance2242();
    output_declaration2243 output_declaration_instance2243();
    output_declaration2244 output_declaration_instance2244();
    output_declaration2245 output_declaration_instance2245();
    output_declaration2246 output_declaration_instance2246();
    output_declaration2247 output_declaration_instance2247();
    output_declaration2248 output_declaration_instance2248();
    output_declaration2249 output_declaration_instance2249();
    output_declaration2250 output_declaration_instance2250();
    output_declaration2251 output_declaration_instance2251();
    output_declaration2252 output_declaration_instance2252();
    output_declaration2253 output_declaration_instance2253();
    output_declaration2254 output_declaration_instance2254();
    output_declaration2255 output_declaration_instance2255();
    output_declaration2256 output_declaration_instance2256();
    output_declaration2257 output_declaration_instance2257();
    output_declaration2258 output_declaration_instance2258();
    output_declaration2259 output_declaration_instance2259();
    output_declaration2260 output_declaration_instance2260();
    output_declaration2261 output_declaration_instance2261();
    output_declaration2262 output_declaration_instance2262();
    output_declaration2263 output_declaration_instance2263();
    output_declaration2264 output_declaration_instance2264();
    output_declaration2265 output_declaration_instance2265();
    output_declaration2266 output_declaration_instance2266();
    output_declaration2267 output_declaration_instance2267();
    output_declaration2268 output_declaration_instance2268();
    output_declaration2269 output_declaration_instance2269();
    output_declaration2270 output_declaration_instance2270();
    output_declaration2271 output_declaration_instance2271();
    output_declaration2272 output_declaration_instance2272();
    output_declaration2273 output_declaration_instance2273();
    output_declaration2274 output_declaration_instance2274();
    output_declaration2275 output_declaration_instance2275();
    output_declaration2276 output_declaration_instance2276();
    output_declaration2277 output_declaration_instance2277();
    output_declaration2278 output_declaration_instance2278();
    output_declaration2279 output_declaration_instance2279();
    output_declaration2280 output_declaration_instance2280();
    output_declaration2281 output_declaration_instance2281();
    output_declaration2282 output_declaration_instance2282();
    output_declaration2283 output_declaration_instance2283();
    output_declaration2284 output_declaration_instance2284();
    output_declaration2285 output_declaration_instance2285();
    output_declaration2286 output_declaration_instance2286();
    output_declaration2287 output_declaration_instance2287();
    output_declaration2288 output_declaration_instance2288();
    output_declaration2289 output_declaration_instance2289();
    output_declaration2290 output_declaration_instance2290();
    output_declaration2291 output_declaration_instance2291();
    output_declaration2292 output_declaration_instance2292();
    output_declaration2293 output_declaration_instance2293();
    output_declaration2294 output_declaration_instance2294();
    output_declaration2295 output_declaration_instance2295();
    output_declaration2296 output_declaration_instance2296();
    output_declaration2297 output_declaration_instance2297();
    output_declaration2298 output_declaration_instance2298();
    output_declaration2299 output_declaration_instance2299();
    output_declaration2300 output_declaration_instance2300();
    output_declaration2301 output_declaration_instance2301();
    output_declaration2302 output_declaration_instance2302();
    output_declaration2303 output_declaration_instance2303();
    output_declaration2304 output_declaration_instance2304();
    output_declaration2305 output_declaration_instance2305();
    output_declaration2306 output_declaration_instance2306();
    output_declaration2307 output_declaration_instance2307();
    output_declaration2308 output_declaration_instance2308();
    output_declaration2309 output_declaration_instance2309();
    output_declaration2310 output_declaration_instance2310();
    output_declaration2311 output_declaration_instance2311();
    output_declaration2312 output_declaration_instance2312();
    output_declaration2313 output_declaration_instance2313();
    output_declaration2314 output_declaration_instance2314();
    output_declaration2315 output_declaration_instance2315();
    output_declaration2316 output_declaration_instance2316();
    output_declaration2317 output_declaration_instance2317();
    output_declaration2318 output_declaration_instance2318();
    output_declaration2319 output_declaration_instance2319();
    output_declaration2320 output_declaration_instance2320();
    output_declaration2321 output_declaration_instance2321();
    output_declaration2322 output_declaration_instance2322();
    output_declaration2323 output_declaration_instance2323();
    output_declaration2324 output_declaration_instance2324();
    output_declaration2325 output_declaration_instance2325();
    output_declaration2326 output_declaration_instance2326();
    output_declaration2327 output_declaration_instance2327();
    output_declaration2328 output_declaration_instance2328();
    output_declaration2329 output_declaration_instance2329();
    output_declaration2330 output_declaration_instance2330();
    output_declaration2331 output_declaration_instance2331();
    output_declaration2332 output_declaration_instance2332();
    output_declaration2333 output_declaration_instance2333();
    output_declaration2334 output_declaration_instance2334();
    output_declaration2335 output_declaration_instance2335();
    output_declaration2336 output_declaration_instance2336();
    output_declaration2337 output_declaration_instance2337();
    output_declaration2338 output_declaration_instance2338();
    output_declaration2339 output_declaration_instance2339();
    output_declaration2340 output_declaration_instance2340();
    output_declaration2341 output_declaration_instance2341();
    output_declaration2342 output_declaration_instance2342();
    output_declaration2343 output_declaration_instance2343();
    output_declaration2344 output_declaration_instance2344();
    output_declaration2345 output_declaration_instance2345();
    output_declaration2346 output_declaration_instance2346();
    output_declaration2347 output_declaration_instance2347();
    output_declaration2348 output_declaration_instance2348();
    output_declaration2349 output_declaration_instance2349();
    output_declaration2350 output_declaration_instance2350();
    output_declaration2351 output_declaration_instance2351();
    output_declaration2352 output_declaration_instance2352();
    output_declaration2353 output_declaration_instance2353();
    output_declaration2354 output_declaration_instance2354();
    output_declaration2355 output_declaration_instance2355();
    output_declaration2356 output_declaration_instance2356();
    output_declaration2357 output_declaration_instance2357();
    output_declaration2358 output_declaration_instance2358();
    output_declaration2359 output_declaration_instance2359();
    output_declaration2360 output_declaration_instance2360();
    output_declaration2361 output_declaration_instance2361();
    output_declaration2362 output_declaration_instance2362();
    output_declaration2363 output_declaration_instance2363();
    output_declaration2364 output_declaration_instance2364();
    output_declaration2365 output_declaration_instance2365();
    output_declaration2366 output_declaration_instance2366();
    output_declaration2367 output_declaration_instance2367();
    output_declaration2368 output_declaration_instance2368();
    output_declaration2369 output_declaration_instance2369();
    output_declaration2370 output_declaration_instance2370();
    output_declaration2371 output_declaration_instance2371();
    output_declaration2372 output_declaration_instance2372();
    output_declaration2373 output_declaration_instance2373();
    output_declaration2374 output_declaration_instance2374();
    output_declaration2375 output_declaration_instance2375();
    output_declaration2376 output_declaration_instance2376();
    output_declaration2377 output_declaration_instance2377();
    output_declaration2378 output_declaration_instance2378();
    output_declaration2379 output_declaration_instance2379();
    output_declaration2380 output_declaration_instance2380();
    output_declaration2381 output_declaration_instance2381();
    output_declaration2382 output_declaration_instance2382();
    output_declaration2383 output_declaration_instance2383();
    output_declaration2384 output_declaration_instance2384();
    output_declaration2385 output_declaration_instance2385();
    output_declaration2386 output_declaration_instance2386();
    output_declaration2387 output_declaration_instance2387();
    output_declaration2388 output_declaration_instance2388();
    output_declaration2389 output_declaration_instance2389();
    output_declaration2390 output_declaration_instance2390();
    output_declaration2391 output_declaration_instance2391();
    output_declaration2392 output_declaration_instance2392();
    output_declaration2393 output_declaration_instance2393();
    output_declaration2394 output_declaration_instance2394();
    output_declaration2395 output_declaration_instance2395();
    output_declaration2396 output_declaration_instance2396();
    output_declaration2397 output_declaration_instance2397();
    output_declaration2398 output_declaration_instance2398();
    output_declaration2399 output_declaration_instance2399();
    output_declaration2400 output_declaration_instance2400();
    output_declaration2401 output_declaration_instance2401();
    output_declaration2402 output_declaration_instance2402();
    output_declaration2403 output_declaration_instance2403();
    output_declaration2404 output_declaration_instance2404();
    output_declaration2405 output_declaration_instance2405();
    output_declaration2406 output_declaration_instance2406();
    output_declaration2407 output_declaration_instance2407();
    output_declaration2408 output_declaration_instance2408();
    output_declaration2409 output_declaration_instance2409();
    output_declaration2410 output_declaration_instance2410();
    output_declaration2411 output_declaration_instance2411();
    output_declaration2412 output_declaration_instance2412();
    output_declaration2413 output_declaration_instance2413();
    output_declaration2414 output_declaration_instance2414();
    output_declaration2415 output_declaration_instance2415();
    output_declaration2416 output_declaration_instance2416();
    output_declaration2417 output_declaration_instance2417();
    output_declaration2418 output_declaration_instance2418();
    output_declaration2419 output_declaration_instance2419();
    output_declaration2420 output_declaration_instance2420();
    output_declaration2421 output_declaration_instance2421();
    output_declaration2422 output_declaration_instance2422();
    output_declaration2423 output_declaration_instance2423();
    output_declaration2424 output_declaration_instance2424();
    output_declaration2425 output_declaration_instance2425();
    output_declaration2426 output_declaration_instance2426();
    output_declaration2427 output_declaration_instance2427();
    output_declaration2428 output_declaration_instance2428();
    output_declaration2429 output_declaration_instance2429();
    output_declaration2430 output_declaration_instance2430();
    output_declaration2431 output_declaration_instance2431();
    output_declaration2432 output_declaration_instance2432();
    output_declaration2433 output_declaration_instance2433();
    output_declaration2434 output_declaration_instance2434();
    output_declaration2435 output_declaration_instance2435();
    output_declaration2436 output_declaration_instance2436();
    output_declaration2437 output_declaration_instance2437();
    output_declaration2438 output_declaration_instance2438();
    output_declaration2439 output_declaration_instance2439();
    output_declaration2440 output_declaration_instance2440();
    output_declaration2441 output_declaration_instance2441();
    output_declaration2442 output_declaration_instance2442();
    output_declaration2443 output_declaration_instance2443();
    output_declaration2444 output_declaration_instance2444();
    output_declaration2445 output_declaration_instance2445();
    output_declaration2446 output_declaration_instance2446();
    output_declaration2447 output_declaration_instance2447();
    output_declaration2448 output_declaration_instance2448();
    output_declaration2449 output_declaration_instance2449();
    output_declaration2450 output_declaration_instance2450();
    output_declaration2451 output_declaration_instance2451();
    output_declaration2452 output_declaration_instance2452();
    output_declaration2453 output_declaration_instance2453();
    output_declaration2454 output_declaration_instance2454();
    output_declaration2455 output_declaration_instance2455();
    output_declaration2456 output_declaration_instance2456();
    output_declaration2457 output_declaration_instance2457();
    output_declaration2458 output_declaration_instance2458();
    output_declaration2459 output_declaration_instance2459();
    output_declaration2460 output_declaration_instance2460();
    output_declaration2461 output_declaration_instance2461();
    output_declaration2462 output_declaration_instance2462();
    output_declaration2463 output_declaration_instance2463();
    output_declaration2464 output_declaration_instance2464();
    output_declaration2465 output_declaration_instance2465();
    output_declaration2466 output_declaration_instance2466();
    output_declaration2467 output_declaration_instance2467();
    output_declaration2468 output_declaration_instance2468();
    output_declaration2469 output_declaration_instance2469();
    output_declaration2470 output_declaration_instance2470();
    output_declaration2471 output_declaration_instance2471();
    output_declaration2472 output_declaration_instance2472();
    output_declaration2473 output_declaration_instance2473();
    output_declaration2474 output_declaration_instance2474();
    output_declaration2475 output_declaration_instance2475();
    output_declaration2476 output_declaration_instance2476();
    output_declaration2477 output_declaration_instance2477();
    output_declaration2478 output_declaration_instance2478();
    output_declaration2479 output_declaration_instance2479();
    output_declaration2480 output_declaration_instance2480();
    output_declaration2481 output_declaration_instance2481();
    output_declaration2482 output_declaration_instance2482();
    output_declaration2483 output_declaration_instance2483();
    output_declaration2484 output_declaration_instance2484();
    output_declaration2485 output_declaration_instance2485();
    output_declaration2486 output_declaration_instance2486();
    output_declaration2487 output_declaration_instance2487();
    output_declaration2488 output_declaration_instance2488();
    output_declaration2489 output_declaration_instance2489();
    output_declaration2490 output_declaration_instance2490();
    output_declaration2491 output_declaration_instance2491();
    output_declaration2492 output_declaration_instance2492();
    output_declaration2493 output_declaration_instance2493();
    output_declaration2494 output_declaration_instance2494();
    output_declaration2495 output_declaration_instance2495();
    output_declaration2496 output_declaration_instance2496();
    output_declaration2497 output_declaration_instance2497();
    output_declaration2498 output_declaration_instance2498();
    output_declaration2499 output_declaration_instance2499();
    output_declaration2500 output_declaration_instance2500();
    output_declaration2501 output_declaration_instance2501();
    output_declaration2502 output_declaration_instance2502();
    output_declaration2503 output_declaration_instance2503();
    output_declaration2504 output_declaration_instance2504();
    output_declaration2505 output_declaration_instance2505();
    output_declaration2506 output_declaration_instance2506();
    output_declaration2507 output_declaration_instance2507();
    output_declaration2508 output_declaration_instance2508();
    output_declaration2509 output_declaration_instance2509();
    output_declaration2510 output_declaration_instance2510();
    output_declaration2511 output_declaration_instance2511();
    output_declaration2512 output_declaration_instance2512();
    output_declaration2513 output_declaration_instance2513();
    output_declaration2514 output_declaration_instance2514();
    output_declaration2515 output_declaration_instance2515();
endmodule
//@
//author : andreib
module output_declaration0( abc,ABCD ); output abc,ABCD;
endmodule
//author : andreib
module output_declaration1( abc,ABCD ); output [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration2( abc,ABCD ); output [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration3( abc,ABCD ); output [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration4( abc,ABCD ); output [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration5( abc,ABCD ); output [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration6( abc,ABCD ); output [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration7( abc,ABCD ); output [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration8( abc,ABCD ); output [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration9( abc,ABCD ); output [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration10( abc,ABCD ); output [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration11( abc,ABCD ); output [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration12( abc,ABCD ); output [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration13( abc,ABCD ); output [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration14( abc,ABCD ); output [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration15( abc,ABCD ); output [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration16( abc,ABCD ); output [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration17( abc,ABCD ); output [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration18( abc,ABCD ); output [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration19( abc,ABCD ); output [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration20( abc,ABCD ); output [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration21( abc,ABCD ); output [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration22( abc,ABCD ); output [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration23( abc,ABCD ); output [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration24( abc,ABCD ); output [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration25( abc,ABCD ); output [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration26( abc,ABCD ); output signed abc,ABCD;
endmodule
//author : andreib
module output_declaration27( abc,ABCD ); output signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration28( abc,ABCD ); output signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration29( abc,ABCD ); output signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration30( abc,ABCD ); output signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration31( abc,ABCD ); output signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration32( abc,ABCD ); output signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration33( abc,ABCD ); output signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration34( abc,ABCD ); output signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration35( abc,ABCD ); output signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration36( abc,ABCD ); output signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration37( abc,ABCD ); output signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration38( abc,ABCD ); output signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration39( abc,ABCD ); output signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration40( abc,ABCD ); output signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration41( abc,ABCD ); output signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration42( abc,ABCD ); output signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration43( abc,ABCD ); output signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration44( abc,ABCD ); output signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration45( abc,ABCD ); output signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration46( abc,ABCD ); output signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration47( abc,ABCD ); output signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration48( abc,ABCD ); output signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration49( abc,ABCD ); output signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration50( abc,ABCD ); output signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration51( abc,ABCD ); output signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration52( abc,ABCD ); output supply0 abc,ABCD;
endmodule
//author : andreib
module output_declaration53( abc,ABCD ); output supply0 [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration54( abc,ABCD ); output supply0 [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration55( abc,ABCD ); output supply0 [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration56( abc,ABCD ); output supply0 [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration57( abc,ABCD ); output supply0 [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration58( abc,ABCD ); output supply0 [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration59( abc,ABCD ); output supply0 [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration60( abc,ABCD ); output supply0 [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration61( abc,ABCD ); output supply0 [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration62( abc,ABCD ); output supply0 [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration63( abc,ABCD ); output supply0 [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration64( abc,ABCD ); output supply0 [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration65( abc,ABCD ); output supply0 [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration66( abc,ABCD ); output supply0 [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration67( abc,ABCD ); output supply0 [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration68( abc,ABCD ); output supply0 [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration69( abc,ABCD ); output supply0 [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration70( abc,ABCD ); output supply0 [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration71( abc,ABCD ); output supply0 [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration72( abc,ABCD ); output supply0 [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration73( abc,ABCD ); output supply0 [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration74( abc,ABCD ); output supply0 [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration75( abc,ABCD ); output supply0 [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration76( abc,ABCD ); output supply0 [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration77( abc,ABCD ); output supply0 [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration78( abc,ABCD ); output supply0 signed abc,ABCD;
endmodule
//author : andreib
module output_declaration79( abc,ABCD ); output supply0 signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration80( abc,ABCD ); output supply0 signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration81( abc,ABCD ); output supply0 signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration82( abc,ABCD ); output supply0 signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration83( abc,ABCD ); output supply0 signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration84( abc,ABCD ); output supply0 signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration85( abc,ABCD ); output supply0 signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration86( abc,ABCD ); output supply0 signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration87( abc,ABCD ); output supply0 signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration88( abc,ABCD ); output supply0 signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration89( abc,ABCD ); output supply0 signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration90( abc,ABCD ); output supply0 signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration91( abc,ABCD ); output supply0 signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration92( abc,ABCD ); output supply0 signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration93( abc,ABCD ); output supply0 signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration94( abc,ABCD ); output supply0 signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration95( abc,ABCD ); output supply0 signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration96( abc,ABCD ); output supply0 signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration97( abc,ABCD ); output supply0 signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration98( abc,ABCD ); output supply0 signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration99( abc,ABCD ); output supply0 signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration100( abc,ABCD ); output supply0 signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration101( abc,ABCD ); output supply0 signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration102( abc,ABCD ); output supply0 signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration103( abc,ABCD ); output supply0 signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration104( abc,ABCD ); output supply1 abc,ABCD;
endmodule
//author : andreib
module output_declaration105( abc,ABCD ); output supply1 [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration106( abc,ABCD ); output supply1 [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration107( abc,ABCD ); output supply1 [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration108( abc,ABCD ); output supply1 [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration109( abc,ABCD ); output supply1 [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration110( abc,ABCD ); output supply1 [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration111( abc,ABCD ); output supply1 [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration112( abc,ABCD ); output supply1 [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration113( abc,ABCD ); output supply1 [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration114( abc,ABCD ); output supply1 [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration115( abc,ABCD ); output supply1 [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration116( abc,ABCD ); output supply1 [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration117( abc,ABCD ); output supply1 [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration118( abc,ABCD ); output supply1 [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration119( abc,ABCD ); output supply1 [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration120( abc,ABCD ); output supply1 [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration121( abc,ABCD ); output supply1 [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration122( abc,ABCD ); output supply1 [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration123( abc,ABCD ); output supply1 [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration124( abc,ABCD ); output supply1 [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration125( abc,ABCD ); output supply1 [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration126( abc,ABCD ); output supply1 [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration127( abc,ABCD ); output supply1 [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration128( abc,ABCD ); output supply1 [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration129( abc,ABCD ); output supply1 [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration130( abc,ABCD ); output supply1 signed abc,ABCD;
endmodule
//author : andreib
module output_declaration131( abc,ABCD ); output supply1 signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration132( abc,ABCD ); output supply1 signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration133( abc,ABCD ); output supply1 signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration134( abc,ABCD ); output supply1 signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration135( abc,ABCD ); output supply1 signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration136( abc,ABCD ); output supply1 signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration137( abc,ABCD ); output supply1 signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration138( abc,ABCD ); output supply1 signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration139( abc,ABCD ); output supply1 signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration140( abc,ABCD ); output supply1 signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration141( abc,ABCD ); output supply1 signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration142( abc,ABCD ); output supply1 signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration143( abc,ABCD ); output supply1 signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration144( abc,ABCD ); output supply1 signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration145( abc,ABCD ); output supply1 signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration146( abc,ABCD ); output supply1 signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration147( abc,ABCD ); output supply1 signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration148( abc,ABCD ); output supply1 signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration149( abc,ABCD ); output supply1 signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration150( abc,ABCD ); output supply1 signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration151( abc,ABCD ); output supply1 signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration152( abc,ABCD ); output supply1 signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration153( abc,ABCD ); output supply1 signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration154( abc,ABCD ); output supply1 signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration155( abc,ABCD ); output supply1 signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration156( abc,ABCD ); output tri abc,ABCD;
endmodule
//author : andreib
module output_declaration157( abc,ABCD ); output tri [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration158( abc,ABCD ); output tri [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration159( abc,ABCD ); output tri [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration160( abc,ABCD ); output tri [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration161( abc,ABCD ); output tri [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration162( abc,ABCD ); output tri [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration163( abc,ABCD ); output tri [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration164( abc,ABCD ); output tri [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration165( abc,ABCD ); output tri [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration166( abc,ABCD ); output tri [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration167( abc,ABCD ); output tri [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration168( abc,ABCD ); output tri [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration169( abc,ABCD ); output tri [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration170( abc,ABCD ); output tri [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration171( abc,ABCD ); output tri [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration172( abc,ABCD ); output tri [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration173( abc,ABCD ); output tri [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration174( abc,ABCD ); output tri [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration175( abc,ABCD ); output tri [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration176( abc,ABCD ); output tri [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration177( abc,ABCD ); output tri [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration178( abc,ABCD ); output tri [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration179( abc,ABCD ); output tri [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration180( abc,ABCD ); output tri [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration181( abc,ABCD ); output tri [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration182( abc,ABCD ); output tri signed abc,ABCD;
endmodule
//author : andreib
module output_declaration183( abc,ABCD ); output tri signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration184( abc,ABCD ); output tri signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration185( abc,ABCD ); output tri signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration186( abc,ABCD ); output tri signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration187( abc,ABCD ); output tri signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration188( abc,ABCD ); output tri signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration189( abc,ABCD ); output tri signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration190( abc,ABCD ); output tri signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration191( abc,ABCD ); output tri signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration192( abc,ABCD ); output tri signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration193( abc,ABCD ); output tri signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration194( abc,ABCD ); output tri signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration195( abc,ABCD ); output tri signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration196( abc,ABCD ); output tri signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration197( abc,ABCD ); output tri signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration198( abc,ABCD ); output tri signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration199( abc,ABCD ); output tri signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration200( abc,ABCD ); output tri signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration201( abc,ABCD ); output tri signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration202( abc,ABCD ); output tri signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration203( abc,ABCD ); output tri signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration204( abc,ABCD ); output tri signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration205( abc,ABCD ); output tri signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration206( abc,ABCD ); output tri signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration207( abc,ABCD ); output tri signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration208( abc,ABCD ); output triand abc,ABCD;
endmodule
//author : andreib
module output_declaration209( abc,ABCD ); output triand [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration210( abc,ABCD ); output triand [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration211( abc,ABCD ); output triand [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration212( abc,ABCD ); output triand [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration213( abc,ABCD ); output triand [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration214( abc,ABCD ); output triand [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration215( abc,ABCD ); output triand [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration216( abc,ABCD ); output triand [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration217( abc,ABCD ); output triand [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration218( abc,ABCD ); output triand [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration219( abc,ABCD ); output triand [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration220( abc,ABCD ); output triand [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration221( abc,ABCD ); output triand [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration222( abc,ABCD ); output triand [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration223( abc,ABCD ); output triand [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration224( abc,ABCD ); output triand [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration225( abc,ABCD ); output triand [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration226( abc,ABCD ); output triand [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration227( abc,ABCD ); output triand [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration228( abc,ABCD ); output triand [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration229( abc,ABCD ); output triand [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration230( abc,ABCD ); output triand [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration231( abc,ABCD ); output triand [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration232( abc,ABCD ); output triand [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration233( abc,ABCD ); output triand [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration234( abc,ABCD ); output triand signed abc,ABCD;
endmodule
//author : andreib
module output_declaration235( abc,ABCD ); output triand signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration236( abc,ABCD ); output triand signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration237( abc,ABCD ); output triand signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration238( abc,ABCD ); output triand signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration239( abc,ABCD ); output triand signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration240( abc,ABCD ); output triand signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration241( abc,ABCD ); output triand signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration242( abc,ABCD ); output triand signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration243( abc,ABCD ); output triand signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration244( abc,ABCD ); output triand signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration245( abc,ABCD ); output triand signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration246( abc,ABCD ); output triand signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration247( abc,ABCD ); output triand signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration248( abc,ABCD ); output triand signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration249( abc,ABCD ); output triand signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration250( abc,ABCD ); output triand signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration251( abc,ABCD ); output triand signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration252( abc,ABCD ); output triand signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration253( abc,ABCD ); output triand signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration254( abc,ABCD ); output triand signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration255( abc,ABCD ); output triand signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration256( abc,ABCD ); output triand signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration257( abc,ABCD ); output triand signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration258( abc,ABCD ); output triand signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration259( abc,ABCD ); output triand signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration260( abc,ABCD ); output trior abc,ABCD;
endmodule
//author : andreib
module output_declaration261( abc,ABCD ); output trior [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration262( abc,ABCD ); output trior [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration263( abc,ABCD ); output trior [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration264( abc,ABCD ); output trior [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration265( abc,ABCD ); output trior [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration266( abc,ABCD ); output trior [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration267( abc,ABCD ); output trior [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration268( abc,ABCD ); output trior [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration269( abc,ABCD ); output trior [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration270( abc,ABCD ); output trior [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration271( abc,ABCD ); output trior [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration272( abc,ABCD ); output trior [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration273( abc,ABCD ); output trior [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration274( abc,ABCD ); output trior [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration275( abc,ABCD ); output trior [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration276( abc,ABCD ); output trior [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration277( abc,ABCD ); output trior [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration278( abc,ABCD ); output trior [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration279( abc,ABCD ); output trior [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration280( abc,ABCD ); output trior [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration281( abc,ABCD ); output trior [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration282( abc,ABCD ); output trior [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration283( abc,ABCD ); output trior [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration284( abc,ABCD ); output trior [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration285( abc,ABCD ); output trior [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration286( abc,ABCD ); output trior signed abc,ABCD;
endmodule
//author : andreib
module output_declaration287( abc,ABCD ); output trior signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration288( abc,ABCD ); output trior signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration289( abc,ABCD ); output trior signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration290( abc,ABCD ); output trior signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration291( abc,ABCD ); output trior signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration292( abc,ABCD ); output trior signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration293( abc,ABCD ); output trior signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration294( abc,ABCD ); output trior signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration295( abc,ABCD ); output trior signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration296( abc,ABCD ); output trior signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration297( abc,ABCD ); output trior signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration298( abc,ABCD ); output trior signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration299( abc,ABCD ); output trior signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration300( abc,ABCD ); output trior signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration301( abc,ABCD ); output trior signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration302( abc,ABCD ); output trior signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration303( abc,ABCD ); output trior signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration304( abc,ABCD ); output trior signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration305( abc,ABCD ); output trior signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration306( abc,ABCD ); output trior signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration307( abc,ABCD ); output trior signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration308( abc,ABCD ); output trior signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration309( abc,ABCD ); output trior signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration310( abc,ABCD ); output trior signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration311( abc,ABCD ); output trior signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration312( abc,ABCD ); output tri0 abc,ABCD;
endmodule
//author : andreib
module output_declaration313( abc,ABCD ); output tri0 [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration314( abc,ABCD ); output tri0 [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration315( abc,ABCD ); output tri0 [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration316( abc,ABCD ); output tri0 [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration317( abc,ABCD ); output tri0 [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration318( abc,ABCD ); output tri0 [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration319( abc,ABCD ); output tri0 [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration320( abc,ABCD ); output tri0 [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration321( abc,ABCD ); output tri0 [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration322( abc,ABCD ); output tri0 [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration323( abc,ABCD ); output tri0 [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration324( abc,ABCD ); output tri0 [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration325( abc,ABCD ); output tri0 [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration326( abc,ABCD ); output tri0 [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration327( abc,ABCD ); output tri0 [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration328( abc,ABCD ); output tri0 [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration329( abc,ABCD ); output tri0 [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration330( abc,ABCD ); output tri0 [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration331( abc,ABCD ); output tri0 [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration332( abc,ABCD ); output tri0 [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration333( abc,ABCD ); output tri0 [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration334( abc,ABCD ); output tri0 [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration335( abc,ABCD ); output tri0 [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration336( abc,ABCD ); output tri0 [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration337( abc,ABCD ); output tri0 [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration338( abc,ABCD ); output tri0 signed abc,ABCD;
endmodule
//author : andreib
module output_declaration339( abc,ABCD ); output tri0 signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration340( abc,ABCD ); output tri0 signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration341( abc,ABCD ); output tri0 signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration342( abc,ABCD ); output tri0 signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration343( abc,ABCD ); output tri0 signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration344( abc,ABCD ); output tri0 signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration345( abc,ABCD ); output tri0 signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration346( abc,ABCD ); output tri0 signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration347( abc,ABCD ); output tri0 signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration348( abc,ABCD ); output tri0 signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration349( abc,ABCD ); output tri0 signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration350( abc,ABCD ); output tri0 signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration351( abc,ABCD ); output tri0 signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration352( abc,ABCD ); output tri0 signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration353( abc,ABCD ); output tri0 signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration354( abc,ABCD ); output tri0 signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration355( abc,ABCD ); output tri0 signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration356( abc,ABCD ); output tri0 signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration357( abc,ABCD ); output tri0 signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration358( abc,ABCD ); output tri0 signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration359( abc,ABCD ); output tri0 signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration360( abc,ABCD ); output tri0 signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration361( abc,ABCD ); output tri0 signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration362( abc,ABCD ); output tri0 signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration363( abc,ABCD ); output tri0 signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration364( abc,ABCD ); output tri1 abc,ABCD;
endmodule
//author : andreib
module output_declaration365( abc,ABCD ); output tri1 [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration366( abc,ABCD ); output tri1 [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration367( abc,ABCD ); output tri1 [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration368( abc,ABCD ); output tri1 [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration369( abc,ABCD ); output tri1 [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration370( abc,ABCD ); output tri1 [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration371( abc,ABCD ); output tri1 [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration372( abc,ABCD ); output tri1 [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration373( abc,ABCD ); output tri1 [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration374( abc,ABCD ); output tri1 [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration375( abc,ABCD ); output tri1 [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration376( abc,ABCD ); output tri1 [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration377( abc,ABCD ); output tri1 [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration378( abc,ABCD ); output tri1 [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration379( abc,ABCD ); output tri1 [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration380( abc,ABCD ); output tri1 [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration381( abc,ABCD ); output tri1 [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration382( abc,ABCD ); output tri1 [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration383( abc,ABCD ); output tri1 [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration384( abc,ABCD ); output tri1 [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration385( abc,ABCD ); output tri1 [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration386( abc,ABCD ); output tri1 [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration387( abc,ABCD ); output tri1 [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration388( abc,ABCD ); output tri1 [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration389( abc,ABCD ); output tri1 [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration390( abc,ABCD ); output tri1 signed abc,ABCD;
endmodule
//author : andreib
module output_declaration391( abc,ABCD ); output tri1 signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration392( abc,ABCD ); output tri1 signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration393( abc,ABCD ); output tri1 signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration394( abc,ABCD ); output tri1 signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration395( abc,ABCD ); output tri1 signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration396( abc,ABCD ); output tri1 signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration397( abc,ABCD ); output tri1 signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration398( abc,ABCD ); output tri1 signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration399( abc,ABCD ); output tri1 signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration400( abc,ABCD ); output tri1 signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration401( abc,ABCD ); output tri1 signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration402( abc,ABCD ); output tri1 signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration403( abc,ABCD ); output tri1 signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration404( abc,ABCD ); output tri1 signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration405( abc,ABCD ); output tri1 signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration406( abc,ABCD ); output tri1 signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration407( abc,ABCD ); output tri1 signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration408( abc,ABCD ); output tri1 signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration409( abc,ABCD ); output tri1 signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration410( abc,ABCD ); output tri1 signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration411( abc,ABCD ); output tri1 signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration412( abc,ABCD ); output tri1 signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration413( abc,ABCD ); output tri1 signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration414( abc,ABCD ); output tri1 signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration415( abc,ABCD ); output tri1 signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration416( abc,ABCD ); output wire abc,ABCD;
endmodule
//author : andreib
module output_declaration417( abc,ABCD ); output wire [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration418( abc,ABCD ); output wire [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration419( abc,ABCD ); output wire [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration420( abc,ABCD ); output wire [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration421( abc,ABCD ); output wire [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration422( abc,ABCD ); output wire [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration423( abc,ABCD ); output wire [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration424( abc,ABCD ); output wire [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration425( abc,ABCD ); output wire [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration426( abc,ABCD ); output wire [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration427( abc,ABCD ); output wire [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration428( abc,ABCD ); output wire [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration429( abc,ABCD ); output wire [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration430( abc,ABCD ); output wire [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration431( abc,ABCD ); output wire [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration432( abc,ABCD ); output wire [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration433( abc,ABCD ); output wire [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration434( abc,ABCD ); output wire [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration435( abc,ABCD ); output wire [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration436( abc,ABCD ); output wire [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration437( abc,ABCD ); output wire [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration438( abc,ABCD ); output wire [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration439( abc,ABCD ); output wire [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration440( abc,ABCD ); output wire [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration441( abc,ABCD ); output wire [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration442( abc,ABCD ); output wire signed abc,ABCD;
endmodule
//author : andreib
module output_declaration443( abc,ABCD ); output wire signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration444( abc,ABCD ); output wire signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration445( abc,ABCD ); output wire signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration446( abc,ABCD ); output wire signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration447( abc,ABCD ); output wire signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration448( abc,ABCD ); output wire signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration449( abc,ABCD ); output wire signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration450( abc,ABCD ); output wire signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration451( abc,ABCD ); output wire signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration452( abc,ABCD ); output wire signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration453( abc,ABCD ); output wire signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration454( abc,ABCD ); output wire signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration455( abc,ABCD ); output wire signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration456( abc,ABCD ); output wire signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration457( abc,ABCD ); output wire signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration458( abc,ABCD ); output wire signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration459( abc,ABCD ); output wire signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration460( abc,ABCD ); output wire signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration461( abc,ABCD ); output wire signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration462( abc,ABCD ); output wire signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration463( abc,ABCD ); output wire signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration464( abc,ABCD ); output wire signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration465( abc,ABCD ); output wire signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration466( abc,ABCD ); output wire signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration467( abc,ABCD ); output wire signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration468( abc,ABCD ); output wand abc,ABCD;
endmodule
//author : andreib
module output_declaration469( abc,ABCD ); output wand [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration470( abc,ABCD ); output wand [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration471( abc,ABCD ); output wand [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration472( abc,ABCD ); output wand [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration473( abc,ABCD ); output wand [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration474( abc,ABCD ); output wand [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration475( abc,ABCD ); output wand [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration476( abc,ABCD ); output wand [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration477( abc,ABCD ); output wand [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration478( abc,ABCD ); output wand [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration479( abc,ABCD ); output wand [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration480( abc,ABCD ); output wand [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration481( abc,ABCD ); output wand [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration482( abc,ABCD ); output wand [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration483( abc,ABCD ); output wand [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration484( abc,ABCD ); output wand [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration485( abc,ABCD ); output wand [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration486( abc,ABCD ); output wand [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration487( abc,ABCD ); output wand [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration488( abc,ABCD ); output wand [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration489( abc,ABCD ); output wand [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration490( abc,ABCD ); output wand [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration491( abc,ABCD ); output wand [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration492( abc,ABCD ); output wand [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration493( abc,ABCD ); output wand [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration494( abc,ABCD ); output wand signed abc,ABCD;
endmodule
//author : andreib
module output_declaration495( abc,ABCD ); output wand signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration496( abc,ABCD ); output wand signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration497( abc,ABCD ); output wand signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration498( abc,ABCD ); output wand signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration499( abc,ABCD ); output wand signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration500( abc,ABCD ); output wand signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration501( abc,ABCD ); output wand signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration502( abc,ABCD ); output wand signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration503( abc,ABCD ); output wand signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration504( abc,ABCD ); output wand signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration505( abc,ABCD ); output wand signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration506( abc,ABCD ); output wand signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration507( abc,ABCD ); output wand signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration508( abc,ABCD ); output wand signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration509( abc,ABCD ); output wand signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration510( abc,ABCD ); output wand signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration511( abc,ABCD ); output wand signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration512( abc,ABCD ); output wand signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration513( abc,ABCD ); output wand signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration514( abc,ABCD ); output wand signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration515( abc,ABCD ); output wand signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration516( abc,ABCD ); output wand signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration517( abc,ABCD ); output wand signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration518( abc,ABCD ); output wand signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration519( abc,ABCD ); output wand signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration520( abc,ABCD ); output wor abc,ABCD;
endmodule
//author : andreib
module output_declaration521( abc,ABCD ); output wor [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration522( abc,ABCD ); output wor [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration523( abc,ABCD ); output wor [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration524( abc,ABCD ); output wor [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration525( abc,ABCD ); output wor [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration526( abc,ABCD ); output wor [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration527( abc,ABCD ); output wor [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration528( abc,ABCD ); output wor [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration529( abc,ABCD ); output wor [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration530( abc,ABCD ); output wor [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration531( abc,ABCD ); output wor [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration532( abc,ABCD ); output wor [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration533( abc,ABCD ); output wor [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration534( abc,ABCD ); output wor [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration535( abc,ABCD ); output wor [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration536( abc,ABCD ); output wor [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration537( abc,ABCD ); output wor [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration538( abc,ABCD ); output wor [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration539( abc,ABCD ); output wor [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration540( abc,ABCD ); output wor [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration541( abc,ABCD ); output wor [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration542( abc,ABCD ); output wor [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration543( abc,ABCD ); output wor [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration544( abc,ABCD ); output wor [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration545( abc,ABCD ); output wor [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration546( abc,ABCD ); output wor signed abc,ABCD;
endmodule
//author : andreib
module output_declaration547( abc,ABCD ); output wor signed [ 2 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration548( abc,ABCD ); output wor signed [ 2 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration549( abc,ABCD ); output wor signed [ 2 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration550( abc,ABCD ); output wor signed [ 2 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration551( abc,ABCD ); output wor signed [ 2 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration552( abc,ABCD ); output wor signed [ +3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration553( abc,ABCD ); output wor signed [ +3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration554( abc,ABCD ); output wor signed [ +3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration555( abc,ABCD ); output wor signed [ +3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration556( abc,ABCD ); output wor signed [ +3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration557( abc,ABCD ); output wor signed [ 2-1 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration558( abc,ABCD ); output wor signed [ 2-1 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration559( abc,ABCD ); output wor signed [ 2-1 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration560( abc,ABCD ); output wor signed [ 2-1 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration561( abc,ABCD ); output wor signed [ 2-1 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration562( abc,ABCD ); output wor signed [ 1?2:3 : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration563( abc,ABCD ); output wor signed [ 1?2:3 : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration564( abc,ABCD ); output wor signed [ 1?2:3 : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration565( abc,ABCD ); output wor signed [ 1?2:3 : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration566( abc,ABCD ); output wor signed [ 1?2:3 : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration567( abc,ABCD ); output wor signed [ "str" : 1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration568( abc,ABCD ); output wor signed [ "str" : +1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration569( abc,ABCD ); output wor signed [ "str" : 2-1 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration570( abc,ABCD ); output wor signed [ "str" : 1?2:3 ] abc,ABCD;
endmodule
//author : andreib
module output_declaration571( abc,ABCD ); output wor signed [ "str" : "str" ] abc,ABCD;
endmodule
//author : andreib
module output_declaration572( xyz,XYZ ); output reg xyz ,XYZ;
endmodule
//author : andreib
module output_declaration573( xyz,XYZ ); output reg xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration574( xyz,XYZ ); output reg xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration575( xyz,XYZ ); output reg xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration576( xyz,XYZ ); output reg xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration577( xyz,XYZ ); output reg xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration578( xyz,XYZ ); output reg xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration579( xyz,XYZ ); output reg xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration580( xyz,XYZ ); output reg xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration581( xyz,XYZ ); output reg xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration582( xyz,XYZ ); output reg xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration583( xyz,XYZ ); output reg xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration584( xyz,XYZ ); output reg xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration585( xyz,XYZ ); output reg xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration586( xyz,XYZ ); output reg xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration587( xyz,XYZ ); output reg xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration588( xyz,XYZ ); output reg xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration589( xyz,XYZ ); output reg xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration590( xyz,XYZ ); output reg xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration591( xyz,XYZ ); output reg xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration592( xyz,XYZ ); output reg xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration593( xyz,XYZ ); output reg xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration594( xyz,XYZ ); output reg xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration595( xyz,XYZ ); output reg xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration596( xyz,XYZ ); output reg xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration597( xyz,XYZ ); output reg xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration598( xyz,XYZ ); output reg xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration599( xyz,XYZ ); output reg xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration600( xyz,XYZ ); output reg xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration601( xyz,XYZ ); output reg xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration602( xyz,XYZ ); output reg xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration603( xyz,XYZ ); output reg xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration604( xyz,XYZ ); output reg xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration605( xyz,XYZ ); output reg xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration606( xyz,XYZ ); output reg xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration607( xyz,XYZ ); output reg xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration608( xyz,XYZ ); output reg [ 2 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration609( xyz,XYZ ); output reg [ 2 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration610( xyz,XYZ ); output reg [ 2 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration611( xyz,XYZ ); output reg [ 2 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration612( xyz,XYZ ); output reg [ 2 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration613( xyz,XYZ ); output reg [ 2 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration614( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration615( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration616( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration617( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration618( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration619( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration620( xyz,XYZ ); output reg [ 2 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration621( xyz,XYZ ); output reg [ 2 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration622( xyz,XYZ ); output reg [ 2 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration623( xyz,XYZ ); output reg [ 2 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration624( xyz,XYZ ); output reg [ 2 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration625( xyz,XYZ ); output reg [ 2 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration626( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration627( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration628( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration629( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration630( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration631( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration632( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration633( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration634( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration635( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration636( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration637( xyz,XYZ ); output reg [ 2 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration638( xyz,XYZ ); output reg [ 2 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration639( xyz,XYZ ); output reg [ 2 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration640( xyz,XYZ ); output reg [ 2 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration641( xyz,XYZ ); output reg [ 2 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration642( xyz,XYZ ); output reg [ 2 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration643( xyz,XYZ ); output reg [ 2 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration644( xyz,XYZ ); output reg [ 2 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration645( xyz,XYZ ); output reg [ 2 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration646( xyz,XYZ ); output reg [ 2 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration647( xyz,XYZ ); output reg [ 2 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration648( xyz,XYZ ); output reg [ 2 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration649( xyz,XYZ ); output reg [ 2 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration650( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration651( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration652( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration653( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration654( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration655( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration656( xyz,XYZ ); output reg [ 2 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration657( xyz,XYZ ); output reg [ 2 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration658( xyz,XYZ ); output reg [ 2 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration659( xyz,XYZ ); output reg [ 2 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration660( xyz,XYZ ); output reg [ 2 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration661( xyz,XYZ ); output reg [ 2 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration662( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration663( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration664( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration665( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration666( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration667( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration668( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration669( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration670( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration671( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration672( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration673( xyz,XYZ ); output reg [ 2 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration674( xyz,XYZ ); output reg [ 2 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration675( xyz,XYZ ); output reg [ 2 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration676( xyz,XYZ ); output reg [ 2 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration677( xyz,XYZ ); output reg [ 2 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration678( xyz,XYZ ); output reg [ 2 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration679( xyz,XYZ ); output reg [ 2 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration680( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration681( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration682( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration683( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration684( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration685( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration686( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration687( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration688( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration689( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration690( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration691( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration692( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration693( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration694( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration695( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration696( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration697( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration698( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration699( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration700( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration701( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration702( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration703( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration704( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration705( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration706( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration707( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration708( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration709( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration710( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration711( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration712( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration713( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration714( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration715( xyz,XYZ ); output reg [ 2 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration716( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration717( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration718( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration719( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration720( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration721( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration722( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration723( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration724( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration725( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration726( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration727( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration728( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration729( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration730( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration731( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration732( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration733( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration734( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration735( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration736( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration737( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration738( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration739( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration740( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration741( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration742( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration743( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration744( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration745( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration746( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration747( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration748( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration749( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration750( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration751( xyz,XYZ ); output reg [ 2 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration752( xyz,XYZ ); output reg [ 2 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration753( xyz,XYZ ); output reg [ 2 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration754( xyz,XYZ ); output reg [ 2 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration755( xyz,XYZ ); output reg [ 2 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration756( xyz,XYZ ); output reg [ 2 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration757( xyz,XYZ ); output reg [ 2 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration758( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration759( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration760( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration761( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration762( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration763( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration764( xyz,XYZ ); output reg [ 2 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration765( xyz,XYZ ); output reg [ 2 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration766( xyz,XYZ ); output reg [ 2 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration767( xyz,XYZ ); output reg [ 2 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration768( xyz,XYZ ); output reg [ 2 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration769( xyz,XYZ ); output reg [ 2 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration770( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration771( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration772( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration773( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration774( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration775( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration776( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration777( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration778( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration779( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration780( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration781( xyz,XYZ ); output reg [ 2 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration782( xyz,XYZ ); output reg [ 2 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration783( xyz,XYZ ); output reg [ 2 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration784( xyz,XYZ ); output reg [ 2 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration785( xyz,XYZ ); output reg [ 2 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration786( xyz,XYZ ); output reg [ 2 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration787( xyz,XYZ ); output reg [ 2 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration788( xyz,XYZ ); output reg [ +3 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration789( xyz,XYZ ); output reg [ +3 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration790( xyz,XYZ ); output reg [ +3 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration791( xyz,XYZ ); output reg [ +3 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration792( xyz,XYZ ); output reg [ +3 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration793( xyz,XYZ ); output reg [ +3 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration794( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration795( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration796( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration797( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration798( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration799( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration800( xyz,XYZ ); output reg [ +3 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration801( xyz,XYZ ); output reg [ +3 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration802( xyz,XYZ ); output reg [ +3 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration803( xyz,XYZ ); output reg [ +3 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration804( xyz,XYZ ); output reg [ +3 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration805( xyz,XYZ ); output reg [ +3 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration806( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration807( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration808( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration809( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration810( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration811( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration812( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration813( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration814( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration815( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration816( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration817( xyz,XYZ ); output reg [ +3 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration818( xyz,XYZ ); output reg [ +3 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration819( xyz,XYZ ); output reg [ +3 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration820( xyz,XYZ ); output reg [ +3 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration821( xyz,XYZ ); output reg [ +3 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration822( xyz,XYZ ); output reg [ +3 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration823( xyz,XYZ ); output reg [ +3 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration824( xyz,XYZ ); output reg [ +3 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration825( xyz,XYZ ); output reg [ +3 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration826( xyz,XYZ ); output reg [ +3 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration827( xyz,XYZ ); output reg [ +3 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration828( xyz,XYZ ); output reg [ +3 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration829( xyz,XYZ ); output reg [ +3 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration830( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration831( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration832( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration833( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration834( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration835( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration836( xyz,XYZ ); output reg [ +3 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration837( xyz,XYZ ); output reg [ +3 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration838( xyz,XYZ ); output reg [ +3 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration839( xyz,XYZ ); output reg [ +3 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration840( xyz,XYZ ); output reg [ +3 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration841( xyz,XYZ ); output reg [ +3 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration842( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration843( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration844( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration845( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration846( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration847( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration848( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration849( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration850( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration851( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration852( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration853( xyz,XYZ ); output reg [ +3 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration854( xyz,XYZ ); output reg [ +3 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration855( xyz,XYZ ); output reg [ +3 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration856( xyz,XYZ ); output reg [ +3 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration857( xyz,XYZ ); output reg [ +3 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration858( xyz,XYZ ); output reg [ +3 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration859( xyz,XYZ ); output reg [ +3 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration860( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration861( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration862( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration863( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration864( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration865( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration866( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration867( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration868( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration869( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration870( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration871( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration872( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration873( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration874( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration875( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration876( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration877( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration878( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration879( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration880( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration881( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration882( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration883( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration884( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration885( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration886( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration887( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration888( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration889( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration890( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration891( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration892( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration893( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration894( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration895( xyz,XYZ ); output reg [ +3 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration896( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration897( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration898( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration899( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration900( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration901( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration902( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration903( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration904( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration905( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration906( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration907( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration908( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration909( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration910( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration911( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration912( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration913( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration914( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration915( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration916( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration917( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration918( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration919( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration920( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration921( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration922( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration923( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration924( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration925( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration926( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration927( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration928( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration929( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration930( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration931( xyz,XYZ ); output reg [ +3 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration932( xyz,XYZ ); output reg [ +3 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration933( xyz,XYZ ); output reg [ +3 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration934( xyz,XYZ ); output reg [ +3 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration935( xyz,XYZ ); output reg [ +3 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration936( xyz,XYZ ); output reg [ +3 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration937( xyz,XYZ ); output reg [ +3 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration938( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration939( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration940( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration941( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration942( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration943( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration944( xyz,XYZ ); output reg [ +3 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration945( xyz,XYZ ); output reg [ +3 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration946( xyz,XYZ ); output reg [ +3 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration947( xyz,XYZ ); output reg [ +3 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration948( xyz,XYZ ); output reg [ +3 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration949( xyz,XYZ ); output reg [ +3 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration950( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration951( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration952( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration953( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration954( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration955( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration956( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration957( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration958( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration959( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration960( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration961( xyz,XYZ ); output reg [ +3 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration962( xyz,XYZ ); output reg [ +3 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration963( xyz,XYZ ); output reg [ +3 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration964( xyz,XYZ ); output reg [ +3 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration965( xyz,XYZ ); output reg [ +3 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration966( xyz,XYZ ); output reg [ +3 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration967( xyz,XYZ ); output reg [ +3 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration968( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration969( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration970( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration971( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration972( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration973( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration974( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration975( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration976( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration977( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration978( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration979( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration980( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration981( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration982( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration983( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration984( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration985( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration986( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration987( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration988( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration989( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration990( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration991( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration992( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration993( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration994( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration995( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration996( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration997( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration998( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration999( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1000( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1001( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1002( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1003( xyz,XYZ ); output reg [ 2-1 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1004( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1005( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1006( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1007( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1008( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1009( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1010( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1011( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1012( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1013( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1014( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1015( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1016( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1017( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1018( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1019( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1020( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1021( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1022( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1023( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1024( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1025( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1026( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1027( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1028( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1029( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1030( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1031( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1032( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1033( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1034( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1035( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1036( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1037( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1038( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1039( xyz,XYZ ); output reg [ 2-1 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1040( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1041( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1042( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1043( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1044( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1045( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1046( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1047( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1048( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1049( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1050( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1051( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1052( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1053( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1054( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1055( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1056( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1057( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1058( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1059( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1060( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1061( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1062( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1063( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1064( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1065( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1066( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1067( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1068( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1069( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1070( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1071( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1072( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1073( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1074( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1075( xyz,XYZ ); output reg [ 2-1 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1076( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1077( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1078( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1079( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1080( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1081( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1082( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1083( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1084( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1085( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1086( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1087( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1088( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1089( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1090( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1091( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1092( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1093( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1094( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1095( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1096( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1097( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1098( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1099( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1100( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1101( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1102( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1103( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1104( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1105( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1106( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1107( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1108( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1109( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1110( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1111( xyz,XYZ ); output reg [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1112( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1113( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1114( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1115( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1116( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1117( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1118( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1119( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1120( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1121( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1122( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1123( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1124( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1125( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1126( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1127( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1128( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1129( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1130( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1131( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1132( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1133( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1134( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1135( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1136( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1137( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1138( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1139( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1140( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1141( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1142( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1143( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1144( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1145( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1146( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1147( xyz,XYZ ); output reg [ 2-1 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1148( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1149( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1150( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1151( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1152( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1153( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1154( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1155( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1156( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1157( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1158( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1159( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1160( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1161( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1162( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1163( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1164( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1165( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1166( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1167( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1168( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1169( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1170( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1171( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1172( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1173( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1174( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1175( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1176( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1177( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1178( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1179( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1180( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1181( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1182( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1183( xyz,XYZ ); output reg [ 1?2:3 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1184( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1185( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1186( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1187( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1188( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1189( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1190( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1191( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1192( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1193( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1194( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1195( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1196( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1197( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1198( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1199( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1200( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1201( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1202( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1203( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1204( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1205( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1206( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1207( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1208( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1209( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1210( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1211( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1212( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1213( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1214( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1215( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1216( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1217( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1218( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1219( xyz,XYZ ); output reg [ 1?2:3 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1220( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1221( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1222( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1223( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1224( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1225( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1226( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1227( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1228( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1229( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1230( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1231( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1232( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1233( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1234( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1235( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1236( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1237( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1238( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1239( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1240( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1241( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1242( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1243( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1244( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1245( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1246( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1247( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1248( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1249( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1250( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1251( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1252( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1253( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1254( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1255( xyz,XYZ ); output reg [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1256( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1257( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1258( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1259( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1260( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1261( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1262( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1263( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1264( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1265( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1266( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1267( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1268( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1269( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1270( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1271( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1272( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1273( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1274( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1275( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1276( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1277( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1278( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1279( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1280( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1281( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1282( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1283( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1284( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1285( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1286( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1287( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1288( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1289( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1290( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1291( xyz,XYZ ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1292( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1293( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1294( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1295( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1296( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1297( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1298( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1299( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1300( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1301( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1302( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1303( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1304( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1305( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1306( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1307( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1308( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1309( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1310( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1311( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1312( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1313( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1314( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1315( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1316( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1317( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1318( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1319( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1320( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1321( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1322( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1323( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1324( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1325( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1326( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1327( xyz,XYZ ); output reg [ 1?2:3 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1328( xyz,XYZ ); output reg [ "str" : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1329( xyz,XYZ ); output reg [ "str" : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1330( xyz,XYZ ); output reg [ "str" : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1331( xyz,XYZ ); output reg [ "str" : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1332( xyz,XYZ ); output reg [ "str" : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1333( xyz,XYZ ); output reg [ "str" : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1334( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1335( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1336( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1337( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1338( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1339( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1340( xyz,XYZ ); output reg [ "str" : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1341( xyz,XYZ ); output reg [ "str" : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1342( xyz,XYZ ); output reg [ "str" : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1343( xyz,XYZ ); output reg [ "str" : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1344( xyz,XYZ ); output reg [ "str" : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1345( xyz,XYZ ); output reg [ "str" : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1346( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1347( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1348( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1349( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1350( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1351( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1352( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1353( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1354( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1355( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1356( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1357( xyz,XYZ ); output reg [ "str" : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1358( xyz,XYZ ); output reg [ "str" : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1359( xyz,XYZ ); output reg [ "str" : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1360( xyz,XYZ ); output reg [ "str" : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1361( xyz,XYZ ); output reg [ "str" : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1362( xyz,XYZ ); output reg [ "str" : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1363( xyz,XYZ ); output reg [ "str" : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1364( xyz,XYZ ); output reg [ "str" : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1365( xyz,XYZ ); output reg [ "str" : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1366( xyz,XYZ ); output reg [ "str" : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1367( xyz,XYZ ); output reg [ "str" : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1368( xyz,XYZ ); output reg [ "str" : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1369( xyz,XYZ ); output reg [ "str" : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1370( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1371( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1372( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1373( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1374( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1375( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1376( xyz,XYZ ); output reg [ "str" : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1377( xyz,XYZ ); output reg [ "str" : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1378( xyz,XYZ ); output reg [ "str" : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1379( xyz,XYZ ); output reg [ "str" : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1380( xyz,XYZ ); output reg [ "str" : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1381( xyz,XYZ ); output reg [ "str" : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1382( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1383( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1384( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1385( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1386( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1387( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1388( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1389( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1390( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1391( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1392( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1393( xyz,XYZ ); output reg [ "str" : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1394( xyz,XYZ ); output reg [ "str" : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1395( xyz,XYZ ); output reg [ "str" : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1396( xyz,XYZ ); output reg [ "str" : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1397( xyz,XYZ ); output reg [ "str" : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1398( xyz,XYZ ); output reg [ "str" : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1399( xyz,XYZ ); output reg [ "str" : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1400( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1401( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1402( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1403( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1404( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1405( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1406( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1407( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1408( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1409( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1410( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1411( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1412( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1413( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1414( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1415( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1416( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1417( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1418( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1419( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1420( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1421( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1422( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1423( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1424( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1425( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1426( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1427( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1428( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1429( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1430( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1431( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1432( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1433( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1434( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1435( xyz,XYZ ); output reg [ "str" : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1436( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1437( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1438( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1439( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1440( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1441( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1442( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1443( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1444( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1445( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1446( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1447( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1448( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1449( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1450( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1451( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1452( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1453( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1454( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1455( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1456( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1457( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1458( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1459( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1460( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1461( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1462( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1463( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1464( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1465( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1466( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1467( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1468( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1469( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1470( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1471( xyz,XYZ ); output reg [ "str" : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1472( xyz,XYZ ); output reg [ "str" : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1473( xyz,XYZ ); output reg [ "str" : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1474( xyz,XYZ ); output reg [ "str" : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1475( xyz,XYZ ); output reg [ "str" : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1476( xyz,XYZ ); output reg [ "str" : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1477( xyz,XYZ ); output reg [ "str" : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1478( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1479( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1480( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1481( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1482( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1483( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1484( xyz,XYZ ); output reg [ "str" : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1485( xyz,XYZ ); output reg [ "str" : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1486( xyz,XYZ ); output reg [ "str" : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1487( xyz,XYZ ); output reg [ "str" : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1488( xyz,XYZ ); output reg [ "str" : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1489( xyz,XYZ ); output reg [ "str" : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1490( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1491( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1492( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1493( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1494( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1495( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1496( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1497( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1498( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1499( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1500( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1501( xyz,XYZ ); output reg [ "str" : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1502( xyz,XYZ ); output reg [ "str" : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1503( xyz,XYZ ); output reg [ "str" : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1504( xyz,XYZ ); output reg [ "str" : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1505( xyz,XYZ ); output reg [ "str" : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1506( xyz,XYZ ); output reg [ "str" : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1507( xyz,XYZ ); output reg [ "str" : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1508( xyz,XYZ ); output reg signed xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1509( xyz,XYZ ); output reg signed xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1510( xyz,XYZ ); output reg signed xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1511( xyz,XYZ ); output reg signed xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1512( xyz,XYZ ); output reg signed xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1513( xyz,XYZ ); output reg signed xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1514( xyz,XYZ ); output reg signed xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1515( xyz,XYZ ); output reg signed xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1516( xyz,XYZ ); output reg signed xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1517( xyz,XYZ ); output reg signed xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1518( xyz,XYZ ); output reg signed xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1519( xyz,XYZ ); output reg signed xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1520( xyz,XYZ ); output reg signed xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1521( xyz,XYZ ); output reg signed xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1522( xyz,XYZ ); output reg signed xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1523( xyz,XYZ ); output reg signed xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1524( xyz,XYZ ); output reg signed xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1525( xyz,XYZ ); output reg signed xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1526( xyz,XYZ ); output reg signed xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1527( xyz,XYZ ); output reg signed xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1528( xyz,XYZ ); output reg signed xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1529( xyz,XYZ ); output reg signed xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1530( xyz,XYZ ); output reg signed xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1531( xyz,XYZ ); output reg signed xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1532( xyz,XYZ ); output reg signed xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1533( xyz,XYZ ); output reg signed xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1534( xyz,XYZ ); output reg signed xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1535( xyz,XYZ ); output reg signed xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1536( xyz,XYZ ); output reg signed xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1537( xyz,XYZ ); output reg signed xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1538( xyz,XYZ ); output reg signed xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1539( xyz,XYZ ); output reg signed xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1540( xyz,XYZ ); output reg signed xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1541( xyz,XYZ ); output reg signed xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1542( xyz,XYZ ); output reg signed xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1543( xyz,XYZ ); output reg signed xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1544( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1545( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1546( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1547( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1548( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1549( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1550( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1551( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1552( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1553( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1554( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1555( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1556( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1557( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1558( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1559( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1560( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1561( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1562( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1563( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1564( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1565( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1566( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1567( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1568( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1569( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1570( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1571( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1572( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1573( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1574( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1575( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1576( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1577( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1578( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1579( xyz,XYZ ); output reg signed [ 2 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1580( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1581( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1582( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1583( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1584( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1585( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1586( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1587( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1588( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1589( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1590( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1591( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1592( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1593( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1594( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1595( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1596( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1597( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1598( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1599( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1600( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1601( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1602( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1603( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1604( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1605( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1606( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1607( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1608( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1609( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1610( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1611( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1612( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1613( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1614( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1615( xyz,XYZ ); output reg signed [ 2 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1616( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1617( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1618( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1619( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1620( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1621( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1622( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1623( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1624( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1625( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1626( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1627( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1628( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1629( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1630( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1631( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1632( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1633( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1634( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1635( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1636( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1637( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1638( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1639( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1640( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1641( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1642( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1643( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1644( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1645( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1646( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1647( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1648( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1649( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1650( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1651( xyz,XYZ ); output reg signed [ 2 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1652( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1653( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1654( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1655( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1656( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1657( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1658( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1659( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1660( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1661( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1662( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1663( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1664( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1665( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1666( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1667( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1668( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1669( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1670( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1671( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1672( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1673( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1674( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1675( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1676( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1677( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1678( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1679( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1680( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1681( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1682( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1683( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1684( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1685( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1686( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1687( xyz,XYZ ); output reg signed [ 2 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1688( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1689( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1690( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1691( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1692( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1693( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1694( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1695( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1696( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1697( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1698( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1699( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1700( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1701( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1702( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1703( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1704( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1705( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1706( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1707( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1708( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1709( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1710( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1711( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1712( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1713( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1714( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1715( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1716( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1717( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1718( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1719( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1720( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1721( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1722( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1723( xyz,XYZ ); output reg signed [ 2 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1724( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1725( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1726( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1727( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1728( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1729( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1730( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1731( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1732( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1733( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1734( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1735( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1736( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1737( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1738( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1739( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1740( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1741( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1742( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1743( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1744( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1745( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1746( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1747( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1748( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1749( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1750( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1751( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1752( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1753( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1754( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1755( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1756( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1757( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1758( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1759( xyz,XYZ ); output reg signed [ +3 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1760( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1761( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1762( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1763( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1764( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1765( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1766( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1767( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1768( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1769( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1770( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1771( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1772( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1773( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1774( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1775( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1776( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1777( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1778( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1779( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1780( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1781( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1782( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1783( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1784( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1785( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1786( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1787( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1788( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1789( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1790( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1791( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1792( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1793( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1794( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1795( xyz,XYZ ); output reg signed [ +3 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1796( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1797( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1798( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1799( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1800( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1801( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1802( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1803( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1804( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1805( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1806( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1807( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1808( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1809( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1810( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1811( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1812( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1813( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1814( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1815( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1816( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1817( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1818( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1819( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1820( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1821( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1822( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1823( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1824( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1825( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1826( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1827( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1828( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1829( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1830( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1831( xyz,XYZ ); output reg signed [ +3 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1832( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1833( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1834( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1835( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1836( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1837( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1838( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1839( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1840( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1841( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1842( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1843( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1844( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1845( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1846( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1847( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1848( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1849( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1850( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1851( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1852( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1853( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1854( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1855( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1856( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1857( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1858( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1859( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1860( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1861( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1862( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1863( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1864( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1865( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1866( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1867( xyz,XYZ ); output reg signed [ +3 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1868( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1869( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1870( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1871( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1872( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1873( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1874( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1875( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1876( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1877( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1878( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1879( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1880( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1881( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1882( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1883( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1884( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1885( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1886( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1887( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1888( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1889( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1890( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1891( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1892( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1893( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1894( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1895( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1896( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1897( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1898( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1899( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1900( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1901( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1902( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1903( xyz,XYZ ); output reg signed [ +3 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1904( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1905( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1906( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1907( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1908( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1909( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1910( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1911( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1912( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1913( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1914( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1915( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1916( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1917( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1918( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1919( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1920( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1921( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1922( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1923( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1924( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1925( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1926( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1927( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1928( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1929( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1930( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1931( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1932( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1933( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1934( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1935( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1936( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1937( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1938( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1939( xyz,XYZ ); output reg signed [ 2-1 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1940( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1941( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1942( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1943( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1944( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1945( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1946( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1947( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1948( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1949( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1950( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1951( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1952( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1953( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1954( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1955( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1956( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1957( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1958( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1959( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1960( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1961( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1962( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1963( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1964( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration1965( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1966( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1967( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1968( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1969( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1970( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration1971( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1972( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1973( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1974( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1975( xyz,XYZ ); output reg signed [ 2-1 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1976( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration1977( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1978( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1979( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1980( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1981( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1982( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration1983( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1984( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1985( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1986( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1987( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1988( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration1989( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1990( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1991( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1992( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1993( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration1994( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration1995( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration1996( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration1997( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration1998( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration1999( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2000( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2001( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2002( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2003( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2004( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2005( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2006( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2007( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2008( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2009( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2010( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2011( xyz,XYZ ); output reg signed [ 2-1 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2012( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2013( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2014( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2015( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2016( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2017( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2018( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2019( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2020( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2021( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2022( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2023( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2024( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2025( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2026( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2027( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2028( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2029( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2030( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2031( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2032( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2033( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2034( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2035( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2036( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2037( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2038( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2039( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2040( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2041( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2042( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2043( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2044( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2045( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2046( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2047( xyz,XYZ ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2048( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2049( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2050( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2051( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2052( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2053( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2054( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2055( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2056( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2057( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2058( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2059( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2060( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2061( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2062( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2063( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2064( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2065( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2066( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2067( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2068( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2069( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2070( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2071( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2072( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2073( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2074( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2075( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2076( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2077( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2078( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2079( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2080( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2081( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2082( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2083( xyz,XYZ ); output reg signed [ 2-1 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2084( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2085( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2086( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2087( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2088( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2089( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2090( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2091( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2092( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2093( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2094( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2095( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2096( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2097( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2098( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2099( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2100( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2101( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2102( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2103( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2104( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2105( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2106( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2107( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2108( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2109( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2110( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2111( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2112( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2113( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2114( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2115( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2116( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2117( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2118( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2119( xyz,XYZ ); output reg signed [ 1?2:3 : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2120( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2121( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2122( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2123( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2124( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2125( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2126( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2127( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2128( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2129( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2130( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2131( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2132( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2133( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2134( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2135( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2136( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2137( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2138( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2139( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2140( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2141( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2142( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2143( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2144( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2145( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2146( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2147( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2148( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2149( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2150( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2151( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2152( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2153( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2154( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2155( xyz,XYZ ); output reg signed [ 1?2:3 : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2156( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2157( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2158( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2159( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2160( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2161( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2162( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2163( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2164( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2165( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2166( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2167( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2168( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2169( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2170( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2171( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2172( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2173( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2174( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2175( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2176( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2177( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2178( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2179( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2180( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2181( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2182( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2183( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2184( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2185( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2186( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2187( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2188( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2189( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2190( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2191( xyz,XYZ ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2192( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2193( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2194( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2195( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2196( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2197( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2198( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2199( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2200( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2201( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2202( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2203( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2204( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2205( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2206( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2207( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2208( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2209( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2210( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2211( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2212( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2213( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2214( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2215( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2216( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2217( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2218( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2219( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2220( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2221( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2222( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2223( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2224( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2225( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2226( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2227( xyz,XYZ ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2228( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2229( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2230( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2231( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2232( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2233( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2234( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2235( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2236( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2237( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2238( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2239( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2240( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2241( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2242( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2243( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2244( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2245( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2246( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2247( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2248( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2249( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2250( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2251( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2252( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2253( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2254( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2255( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2256( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2257( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2258( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2259( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2260( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2261( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2262( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2263( xyz,XYZ ); output reg signed [ 1?2:3 : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2264( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2265( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2266( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2267( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2268( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2269( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2270( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2271( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2272( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2273( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2274( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2275( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2276( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2277( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2278( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2279( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2280( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2281( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2282( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2283( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2284( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2285( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2286( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2287( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2288( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2289( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2290( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2291( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2292( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2293( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2294( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2295( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2296( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2297( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2298( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2299( xyz,XYZ ); output reg signed [ "str" : 1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2300( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2301( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2302( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2303( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2304( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2305( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2306( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2307( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2308( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2309( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2310( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2311( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2312( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2313( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2314( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2315( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2316( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2317( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2318( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2319( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2320( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2321( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2322( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2323( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2324( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2325( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2326( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2327( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2328( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2329( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2330( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2331( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2332( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2333( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2334( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2335( xyz,XYZ ); output reg signed [ "str" : +1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2336( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2337( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2338( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2339( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2340( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2341( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2342( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2343( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2344( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2345( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2346( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2347( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2348( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2349( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2350( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2351( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2352( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2353( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2354( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2355( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2356( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2357( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2358( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2359( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2360( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2361( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2362( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2363( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2364( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2365( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2366( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2367( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2368( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2369( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2370( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2371( xyz,XYZ ); output reg signed [ "str" : 2-1 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2372( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2373( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2374( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2375( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2376( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2377( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2378( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2379( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2380( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2381( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2382( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2383( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2384( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2385( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2386( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2387( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2388( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2389( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2390( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2391( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2392( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2393( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2394( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2395( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2396( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2397( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2398( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2399( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2400( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2401( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2402( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2403( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2404( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2405( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2406( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2407( xyz,XYZ ); output reg signed [ "str" : 1?2:3 ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2408( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2409( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2410( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2411( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2412( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2413( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2414( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2415( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2416( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2417( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2418( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2419( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2420( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2421( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2422( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2423( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2424( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2425( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2426( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2427( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2428( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2429( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2430( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2431( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2432( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2433( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2434( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2435( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2436( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2437( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2438( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2439( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2440( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2441( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2442( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2443( xyz,XYZ ); output reg signed [ "str" : "str" ] xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2444( xyz,XYZ ); output integer xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2445( xyz,XYZ ); output integer xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2446( xyz,XYZ ); output integer xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2447( xyz,XYZ ); output integer xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2448( xyz,XYZ ); output integer xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2449( xyz,XYZ ); output integer xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2450( xyz,XYZ ); output integer xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2451( xyz,XYZ ); output integer xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2452( xyz,XYZ ); output integer xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2453( xyz,XYZ ); output integer xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2454( xyz,XYZ ); output integer xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2455( xyz,XYZ ); output integer xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2456( xyz,XYZ ); output integer xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2457( xyz,XYZ ); output integer xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2458( xyz,XYZ ); output integer xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2459( xyz,XYZ ); output integer xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2460( xyz,XYZ ); output integer xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2461( xyz,XYZ ); output integer xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2462( xyz,XYZ ); output integer xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2463( xyz,XYZ ); output integer xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2464( xyz,XYZ ); output integer xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2465( xyz,XYZ ); output integer xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2466( xyz,XYZ ); output integer xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2467( xyz,XYZ ); output integer xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2468( xyz,XYZ ); output integer xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2469( xyz,XYZ ); output integer xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2470( xyz,XYZ ); output integer xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2471( xyz,XYZ ); output integer xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2472( xyz,XYZ ); output integer xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2473( xyz,XYZ ); output integer xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2474( xyz,XYZ ); output integer xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2475( xyz,XYZ ); output integer xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2476( xyz,XYZ ); output integer xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2477( xyz,XYZ ); output integer xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2478( xyz,XYZ ); output integer xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2479( xyz,XYZ ); output integer xyz = "str" ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2480( xyz,XYZ ); output time xyz ,XYZ;
endmodule
//author : andreib
module output_declaration2481( xyz,XYZ ); output time xyz ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2482( xyz,XYZ ); output time xyz ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2483( xyz,XYZ ); output time xyz ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2484( xyz,XYZ ); output time xyz ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2485( xyz,XYZ ); output time xyz ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2486( xyz,XYZ ); output time xyz = 2 ,XYZ;
endmodule
//author : andreib
module output_declaration2487( xyz,XYZ ); output time xyz = 2 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2488( xyz,XYZ ); output time xyz = 2 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2489( xyz,XYZ ); output time xyz = 2 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2490( xyz,XYZ ); output time xyz = 2 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2491( xyz,XYZ ); output time xyz = 2 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2492( xyz,XYZ ); output time xyz = +3 ,XYZ;
endmodule
//author : andreib
module output_declaration2493( xyz,XYZ ); output time xyz = +3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2494( xyz,XYZ ); output time xyz = +3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2495( xyz,XYZ ); output time xyz = +3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2496( xyz,XYZ ); output time xyz = +3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2497( xyz,XYZ ); output time xyz = +3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2498( xyz,XYZ ); output time xyz = 2-1 ,XYZ;
endmodule
//author : andreib
module output_declaration2499( xyz,XYZ ); output time xyz = 2-1 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2500( xyz,XYZ ); output time xyz = 2-1 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2501( xyz,XYZ ); output time xyz = 2-1 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2502( xyz,XYZ ); output time xyz = 2-1 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2503( xyz,XYZ ); output time xyz = 2-1 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2504( xyz,XYZ ); output time xyz = 1?2:3 ,XYZ;
endmodule
//author : andreib
module output_declaration2505( xyz,XYZ ); output time xyz = 1?2:3 ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2506( xyz,XYZ ); output time xyz = 1?2:3 ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2507( xyz,XYZ ); output time xyz = 1?2:3 ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2508( xyz,XYZ ); output time xyz = 1?2:3 ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2509( xyz,XYZ ); output time xyz = 1?2:3 ,XYZ = "str";
endmodule
//author : andreib
module output_declaration2510( xyz,XYZ ); output time xyz = "str" ,XYZ;
endmodule
//author : andreib
module output_declaration2511( xyz,XYZ ); output time xyz = "str" ,XYZ = 1;
endmodule
//author : andreib
module output_declaration2512( xyz,XYZ ); output time xyz = "str" ,XYZ = +1;
endmodule
//author : andreib
module output_declaration2513( xyz,XYZ ); output time xyz = "str" ,XYZ = 2-1;
endmodule
//author : andreib
module output_declaration2514( xyz,XYZ ); output time xyz = "str" ,XYZ = 1?2:3;
endmodule
//author : andreib
module output_declaration2515( xyz,XYZ ); output time xyz = "str" ,XYZ = "str";
endmodule
