// Test type: blocking_assignment - expression
// Vparser rule name:
// Author: andreib
module blocking_assignment1;
reg a;
initial a=1'b1;
endmodule
