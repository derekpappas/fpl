//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : msi_fabric_if.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module msi_fabric_if(lbdummy2,
                     fab_addbus80,
                     fab_dropbus80);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 45
  output lbdummy2;
  output [79:0] fab_addbus80;
  output [79:0] fab_dropbus80;
  `include "msi_fabric_if.logic.v"
endmodule

