// Test type: case_statement - casex - default null
// Vparser rule name:
// Author: andreib
module case_statement87;
reg a;
initial casex(a)
	default ;
	endcase
endmodule
