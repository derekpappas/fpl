//st1.vh