u1.vhd
top4.vhd
