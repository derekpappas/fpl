`include "defines.v"

module t0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 135
  input [1 - 1:0] ar_sa0_s10;
  s0 s0(.ar_sa0_s10(ar_sa0_s10));
  `include "t0.logic.vh"
endmodule

