u3.vhd
