// Test type: net_assignment - binary operator, 2 attribute instances
// Vparser rule name:
// Author: andreib
module netasign7;
wire a,b,c,d,e;
assign a=b/(*c, d*)e;
endmodule
