`include "defines.v"

module i1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 232
  output [1 - 1:0] ar_sa0_s10;
  h1 h10(.ar_sa0_s10(ar_sa0_s10));
  `include "i1.logic.vh"
endmodule

