// Test type: Continuous assignment - st0, pl1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous106;
wire a;
assign (strong0, pull1) a=1'b1;
endmodule
