`include "defines.v"

module a(p1);
// Location of source csl unit: file name = conn_pattern_ss.csl line number = 4
  input [8 - 1:0] p1;
  `include "a.logic.v"
endmodule

