//test type : module_or_generate_item ::= parameter_declaration
//vparser rule name : 
//author : Codrin
module test_0560;
 (* start = 1, stop *)
 parameter s = 4'b1011, t = 2;
endmodule
