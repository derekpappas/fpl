//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : eth_rx.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module eth_rx();
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 41
  `include "eth_rx.logic.v"
endmodule

