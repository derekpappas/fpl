module b(i);
    wire y;
    input i;
    assign a.x = i;
endmodule