// Test type: initial statement - blocking_assignment - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon1;
reg [7:0]a;
initial a=2;
endmodule
