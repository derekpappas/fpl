//test type : function_port_list ::= input_declaration
//vparser rule name : 
//author : Codrin
module test_0410;
 function [7:0] pow(
  (* width = 8, size *) input nr,
  (* test *) input s);
  pow = 8'b1;
 endfunction
endmodule
