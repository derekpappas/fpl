-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./top1_cslc_generated/code/vhdl/u.vhd
-- FILE GENERATED ON : Sun May 17 09:05:27 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u\ is
  port(\sss_p_p1\ : in csl_bit;
       \sss_p_p2\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \sss_p_p3\ : out csl_bit_vector(10#32# - 10#1# downto 10#0#));
begin
end entity;

architecture \u_logic\ of \u\ is
begin
end architecture;

