`celldefine
module x;
endmodule
`endcelldefine
`celldefine
module y;
endmodule
`resetall
`celldefine
module z;
endmodule
