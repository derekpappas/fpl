`include "defines.v"

module a1(s10);
// Location of source csl unit: file name = temp.csl line number = 182
  output s10;
  `include "a1.logic.vh"
endmodule

