// Test type: Binary Numbers - with z digits and ? digit
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=5'b011z?;
endmodule
