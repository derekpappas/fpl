fifo_port32_in.vhd
loopback32_agent.vhd
fifo_port32_out.vhd
acc.vhd
dp_fp32_gasket.vhd
agent_long_reach.vhd
agent_cluster2.vhd
