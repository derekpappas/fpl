module z(a,c);
  input a;
  output c;
endmodule
module b;
wire y;
wire m;
  z z0(y,m);
endmodule

//module a();
//    b bo();
//endmodule
//module b();
//    a a0();
//endmodule

//module c(m,n);
//    input m;
//    output n;
//endmodule
//module d();
//    c c0();
//endmodule

//module e();
//    wire f,k;
//    z zo();//modul z nedeclarat
//endmodule

//module f();
//    input o, p;
//endmodule


