module mymodule;

  `include "../legal/unconnected_drive05.v"

reg w;
`nounconnected_drive
endmodule
