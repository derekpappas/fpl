//this is a celldefine legal test
module mod;
endmodule
`celldefine/***///sa
