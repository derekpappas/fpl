`include "defines.v"

module h0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 47
  input [1 - 1:0] ar_sa0_s10;
  g0 g0(.ar_sa0_s10(ar_sa0_s10));
  `include "h0.logic.vh"
endmodule

