// Test type: Decimal Numbers - underscore within value
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'd2___9;
endmodule
