`include "defines.v"

module msf();
// Location of source csl unit: file name = IPX2400.csl line number = 74
  `include "msf.logic.v"
endmodule

