-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./msi_rx_cslc_generated/code/vhdl/sfd_trans.vhd
-- FILE GENERATED ON : Tue Jun 17 01:23:46 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity \sfd_trans\ is
end entity;

architecture \sfd_trans_logic\ of \sfd_trans\ is
end architecture;

