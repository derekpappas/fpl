// Test type: Octal Numbers - underscore within size
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=1_2'o1234;
endmodule
