/****/`unconnected_drive pull0
module x;
endmodule
`unconnected_drive pull1
module xx;
endmodule
`unconnected_drive pull0
module xxx;
endmodule
`nounconnected_drive

