-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./b_cslc_generated/code/vhdl/a.vhd
-- FILE GENERATED ON : Mon Feb 16 21:37:22 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \a\ is
  port(\ifc10_x\ : in csl_bit;
       \ifc10_y\ : out csl_bit);
begin
end entity;

architecture \a_logic\ of \a\ is
begin
end architecture;

