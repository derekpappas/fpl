module top();
 wire m,n;
 a a0(.x(m));
 b b0(.y(n));
endmodule
