//test type : module_or_generate_item ::= module_instantiation
//vparser rule name : 
//author : Codrin
module test_0340;
 (* flatten = 1, test = 0, exit *) a a0();
endmodule

module a;
endmodule
