`include "defines.v"

module top();
// Location of source csl unit: file name = set_enum_item_to_field.csl line number = 38
  `include "top.logic.v"
endmodule

