//test type : operator_+ hierarchical_identifier
//vparser rule name : 
//author : Bogdan Mereghea
module unary_operator4;
    wire a, b;
    assign a = +b;
endmodule
