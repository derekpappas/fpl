// Test type: Octal Numbers - 2 numbers, upper case base
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=6'O57;
endmodule
