    `unconnected_drive    pull0         
module x;
endmodule
`resetall
`celldefine
`unconnected_drive    pull1  //
`timescale 10ms/1us
module y;
endmodule
`nounconnected_drive

