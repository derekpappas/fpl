module testbench_output_declaration;
    output_declaration0 output_declaration_instance0();
    output_declaration1 output_declaration_instance1();
    output_declaration2 output_declaration_instance2();
    output_declaration3 output_declaration_instance3();
    output_declaration4 output_declaration_instance4();
    output_declaration5 output_declaration_instance5();
    output_declaration6 output_declaration_instance6();
    output_declaration7 output_declaration_instance7();
    output_declaration8 output_declaration_instance8();
    output_declaration9 output_declaration_instance9();
    output_declaration10 output_declaration_instance10();
    output_declaration11 output_declaration_instance11();
    output_declaration12 output_declaration_instance12();
    output_declaration13 output_declaration_instance13();
    output_declaration14 output_declaration_instance14();
    output_declaration15 output_declaration_instance15();
    output_declaration16 output_declaration_instance16();
    output_declaration17 output_declaration_instance17();
    output_declaration18 output_declaration_instance18();
    output_declaration19 output_declaration_instance19();
    output_declaration20 output_declaration_instance20();
    output_declaration21 output_declaration_instance21();
    output_declaration22 output_declaration_instance22();
    output_declaration23 output_declaration_instance23();
    output_declaration24 output_declaration_instance24();
    output_declaration25 output_declaration_instance25();
    output_declaration26 output_declaration_instance26();
    output_declaration27 output_declaration_instance27();
    output_declaration28 output_declaration_instance28();
    output_declaration29 output_declaration_instance29();
    output_declaration30 output_declaration_instance30();
    output_declaration31 output_declaration_instance31();
    output_declaration32 output_declaration_instance32();
    output_declaration33 output_declaration_instance33();
    output_declaration34 output_declaration_instance34();
    output_declaration35 output_declaration_instance35();
    output_declaration36 output_declaration_instance36();
    output_declaration37 output_declaration_instance37();
    output_declaration38 output_declaration_instance38();
    output_declaration39 output_declaration_instance39();
    output_declaration40 output_declaration_instance40();
    output_declaration41 output_declaration_instance41();
    output_declaration42 output_declaration_instance42();
    output_declaration43 output_declaration_instance43();
    output_declaration44 output_declaration_instance44();
    output_declaration45 output_declaration_instance45();
    output_declaration46 output_declaration_instance46();
    output_declaration47 output_declaration_instance47();
    output_declaration48 output_declaration_instance48();
    output_declaration49 output_declaration_instance49();
    output_declaration50 output_declaration_instance50();
    output_declaration51 output_declaration_instance51();
    output_declaration52 output_declaration_instance52();
    output_declaration53 output_declaration_instance53();
    output_declaration54 output_declaration_instance54();
    output_declaration55 output_declaration_instance55();
    output_declaration56 output_declaration_instance56();
    output_declaration57 output_declaration_instance57();
    output_declaration58 output_declaration_instance58();
    output_declaration59 output_declaration_instance59();
    output_declaration60 output_declaration_instance60();
    output_declaration61 output_declaration_instance61();
    output_declaration62 output_declaration_instance62();
    output_declaration63 output_declaration_instance63();
    output_declaration64 output_declaration_instance64();
    output_declaration65 output_declaration_instance65();
    output_declaration66 output_declaration_instance66();
    output_declaration67 output_declaration_instance67();
    output_declaration68 output_declaration_instance68();
    output_declaration69 output_declaration_instance69();
    output_declaration70 output_declaration_instance70();
    output_declaration71 output_declaration_instance71();
    output_declaration72 output_declaration_instance72();
    output_declaration73 output_declaration_instance73();
    output_declaration74 output_declaration_instance74();
    output_declaration75 output_declaration_instance75();
    output_declaration76 output_declaration_instance76();
    output_declaration77 output_declaration_instance77();
    output_declaration78 output_declaration_instance78();
    output_declaration79 output_declaration_instance79();
    output_declaration80 output_declaration_instance80();
    output_declaration81 output_declaration_instance81();
    output_declaration82 output_declaration_instance82();
    output_declaration83 output_declaration_instance83();
    output_declaration84 output_declaration_instance84();
    output_declaration85 output_declaration_instance85();
    output_declaration86 output_declaration_instance86();
    output_declaration87 output_declaration_instance87();
    output_declaration88 output_declaration_instance88();
    output_declaration89 output_declaration_instance89();
    output_declaration90 output_declaration_instance90();
    output_declaration91 output_declaration_instance91();
    output_declaration92 output_declaration_instance92();
    output_declaration93 output_declaration_instance93();
    output_declaration94 output_declaration_instance94();
    output_declaration95 output_declaration_instance95();
    output_declaration96 output_declaration_instance96();
    output_declaration97 output_declaration_instance97();
    output_declaration98 output_declaration_instance98();
    output_declaration99 output_declaration_instance99();
    output_declaration100 output_declaration_instance100();
    output_declaration101 output_declaration_instance101();
    output_declaration102 output_declaration_instance102();
    output_declaration103 output_declaration_instance103();
    output_declaration104 output_declaration_instance104();
    output_declaration105 output_declaration_instance105();
    output_declaration106 output_declaration_instance106();
    output_declaration107 output_declaration_instance107();
    output_declaration108 output_declaration_instance108();
    output_declaration109 output_declaration_instance109();
    output_declaration110 output_declaration_instance110();
    output_declaration111 output_declaration_instance111();
    output_declaration112 output_declaration_instance112();
    output_declaration113 output_declaration_instance113();
    output_declaration114 output_declaration_instance114();
    output_declaration115 output_declaration_instance115();
    output_declaration116 output_declaration_instance116();
    output_declaration117 output_declaration_instance117();
    output_declaration118 output_declaration_instance118();
    output_declaration119 output_declaration_instance119();
    output_declaration120 output_declaration_instance120();
    output_declaration121 output_declaration_instance121();
    output_declaration122 output_declaration_instance122();
    output_declaration123 output_declaration_instance123();
    output_declaration124 output_declaration_instance124();
    output_declaration125 output_declaration_instance125();
    output_declaration126 output_declaration_instance126();
    output_declaration127 output_declaration_instance127();
    output_declaration128 output_declaration_instance128();
    output_declaration129 output_declaration_instance129();
    output_declaration130 output_declaration_instance130();
    output_declaration131 output_declaration_instance131();
    output_declaration132 output_declaration_instance132();
    output_declaration133 output_declaration_instance133();
    output_declaration134 output_declaration_instance134();
    output_declaration135 output_declaration_instance135();
    output_declaration136 output_declaration_instance136();
    output_declaration137 output_declaration_instance137();
    output_declaration138 output_declaration_instance138();
    output_declaration139 output_declaration_instance139();
    output_declaration140 output_declaration_instance140();
    output_declaration141 output_declaration_instance141();
    output_declaration142 output_declaration_instance142();
    output_declaration143 output_declaration_instance143();
    output_declaration144 output_declaration_instance144();
    output_declaration145 output_declaration_instance145();
    output_declaration146 output_declaration_instance146();
    output_declaration147 output_declaration_instance147();
    output_declaration148 output_declaration_instance148();
    output_declaration149 output_declaration_instance149();
    output_declaration150 output_declaration_instance150();
    output_declaration151 output_declaration_instance151();
    output_declaration152 output_declaration_instance152();
    output_declaration153 output_declaration_instance153();
    output_declaration154 output_declaration_instance154();
    output_declaration155 output_declaration_instance155();
    output_declaration156 output_declaration_instance156();
    output_declaration157 output_declaration_instance157();
    output_declaration158 output_declaration_instance158();
    output_declaration159 output_declaration_instance159();
    output_declaration160 output_declaration_instance160();
    output_declaration161 output_declaration_instance161();
    output_declaration162 output_declaration_instance162();
    output_declaration163 output_declaration_instance163();
    output_declaration164 output_declaration_instance164();
    output_declaration165 output_declaration_instance165();
    output_declaration166 output_declaration_instance166();
    output_declaration167 output_declaration_instance167();
    output_declaration168 output_declaration_instance168();
    output_declaration169 output_declaration_instance169();
    output_declaration170 output_declaration_instance170();
    output_declaration171 output_declaration_instance171();
    output_declaration172 output_declaration_instance172();
    output_declaration173 output_declaration_instance173();
    output_declaration174 output_declaration_instance174();
    output_declaration175 output_declaration_instance175();
    output_declaration176 output_declaration_instance176();
    output_declaration177 output_declaration_instance177();
    output_declaration178 output_declaration_instance178();
    output_declaration179 output_declaration_instance179();
    output_declaration180 output_declaration_instance180();
    output_declaration181 output_declaration_instance181();
    output_declaration182 output_declaration_instance182();
    output_declaration183 output_declaration_instance183();
    output_declaration184 output_declaration_instance184();
    output_declaration185 output_declaration_instance185();
    output_declaration186 output_declaration_instance186();
    output_declaration187 output_declaration_instance187();
    output_declaration188 output_declaration_instance188();
    output_declaration189 output_declaration_instance189();
    output_declaration190 output_declaration_instance190();
    output_declaration191 output_declaration_instance191();
    output_declaration192 output_declaration_instance192();
    output_declaration193 output_declaration_instance193();
    output_declaration194 output_declaration_instance194();
    output_declaration195 output_declaration_instance195();
    output_declaration196 output_declaration_instance196();
    output_declaration197 output_declaration_instance197();
    output_declaration198 output_declaration_instance198();
    output_declaration199 output_declaration_instance199();
    output_declaration200 output_declaration_instance200();
    output_declaration201 output_declaration_instance201();
    output_declaration202 output_declaration_instance202();
    output_declaration203 output_declaration_instance203();
    output_declaration204 output_declaration_instance204();
    output_declaration205 output_declaration_instance205();
    output_declaration206 output_declaration_instance206();
    output_declaration207 output_declaration_instance207();
    output_declaration208 output_declaration_instance208();
    output_declaration209 output_declaration_instance209();
    output_declaration210 output_declaration_instance210();
    output_declaration211 output_declaration_instance211();
    output_declaration212 output_declaration_instance212();
    output_declaration213 output_declaration_instance213();
    output_declaration214 output_declaration_instance214();
    output_declaration215 output_declaration_instance215();
    output_declaration216 output_declaration_instance216();
    output_declaration217 output_declaration_instance217();
    output_declaration218 output_declaration_instance218();
    output_declaration219 output_declaration_instance219();
    output_declaration220 output_declaration_instance220();
    output_declaration221 output_declaration_instance221();
    output_declaration222 output_declaration_instance222();
    output_declaration223 output_declaration_instance223();
    output_declaration224 output_declaration_instance224();
    output_declaration225 output_declaration_instance225();
    output_declaration226 output_declaration_instance226();
    output_declaration227 output_declaration_instance227();
    output_declaration228 output_declaration_instance228();
    output_declaration229 output_declaration_instance229();
    output_declaration230 output_declaration_instance230();
    output_declaration231 output_declaration_instance231();
    output_declaration232 output_declaration_instance232();
    output_declaration233 output_declaration_instance233();
    output_declaration234 output_declaration_instance234();
    output_declaration235 output_declaration_instance235();
    output_declaration236 output_declaration_instance236();
    output_declaration237 output_declaration_instance237();
    output_declaration238 output_declaration_instance238();
    output_declaration239 output_declaration_instance239();
    output_declaration240 output_declaration_instance240();
    output_declaration241 output_declaration_instance241();
    output_declaration242 output_declaration_instance242();
    output_declaration243 output_declaration_instance243();
    output_declaration244 output_declaration_instance244();
    output_declaration245 output_declaration_instance245();
    output_declaration246 output_declaration_instance246();
    output_declaration247 output_declaration_instance247();
    output_declaration248 output_declaration_instance248();
    output_declaration249 output_declaration_instance249();
    output_declaration250 output_declaration_instance250();
    output_declaration251 output_declaration_instance251();
    output_declaration252 output_declaration_instance252();
    output_declaration253 output_declaration_instance253();
    output_declaration254 output_declaration_instance254();
    output_declaration255 output_declaration_instance255();
    output_declaration256 output_declaration_instance256();
    output_declaration257 output_declaration_instance257();
    output_declaration258 output_declaration_instance258();
    output_declaration259 output_declaration_instance259();
    output_declaration260 output_declaration_instance260();
    output_declaration261 output_declaration_instance261();
    output_declaration262 output_declaration_instance262();
    output_declaration263 output_declaration_instance263();
    output_declaration264 output_declaration_instance264();
    output_declaration265 output_declaration_instance265();
    output_declaration266 output_declaration_instance266();
    output_declaration267 output_declaration_instance267();
    output_declaration268 output_declaration_instance268();
    output_declaration269 output_declaration_instance269();
    output_declaration270 output_declaration_instance270();
    output_declaration271 output_declaration_instance271();
    output_declaration272 output_declaration_instance272();
    output_declaration273 output_declaration_instance273();
    output_declaration274 output_declaration_instance274();
    output_declaration275 output_declaration_instance275();
    output_declaration276 output_declaration_instance276();
    output_declaration277 output_declaration_instance277();
    output_declaration278 output_declaration_instance278();
    output_declaration279 output_declaration_instance279();
    output_declaration280 output_declaration_instance280();
    output_declaration281 output_declaration_instance281();
    output_declaration282 output_declaration_instance282();
    output_declaration283 output_declaration_instance283();
    output_declaration284 output_declaration_instance284();
    output_declaration285 output_declaration_instance285();
    output_declaration286 output_declaration_instance286();
    output_declaration287 output_declaration_instance287();
    output_declaration288 output_declaration_instance288();
    output_declaration289 output_declaration_instance289();
    output_declaration290 output_declaration_instance290();
    output_declaration291 output_declaration_instance291();
    output_declaration292 output_declaration_instance292();
    output_declaration293 output_declaration_instance293();
    output_declaration294 output_declaration_instance294();
    output_declaration295 output_declaration_instance295();
    output_declaration296 output_declaration_instance296();
    output_declaration297 output_declaration_instance297();
    output_declaration298 output_declaration_instance298();
    output_declaration299 output_declaration_instance299();
    output_declaration300 output_declaration_instance300();
    output_declaration301 output_declaration_instance301();
    output_declaration302 output_declaration_instance302();
    output_declaration303 output_declaration_instance303();
    output_declaration304 output_declaration_instance304();
    output_declaration305 output_declaration_instance305();
    output_declaration306 output_declaration_instance306();
    output_declaration307 output_declaration_instance307();
    output_declaration308 output_declaration_instance308();
    output_declaration309 output_declaration_instance309();
    output_declaration310 output_declaration_instance310();
    output_declaration311 output_declaration_instance311();
    output_declaration312 output_declaration_instance312();
    output_declaration313 output_declaration_instance313();
    output_declaration314 output_declaration_instance314();
    output_declaration315 output_declaration_instance315();
    output_declaration316 output_declaration_instance316();
    output_declaration317 output_declaration_instance317();
    output_declaration318 output_declaration_instance318();
    output_declaration319 output_declaration_instance319();
    output_declaration320 output_declaration_instance320();
    output_declaration321 output_declaration_instance321();
    output_declaration322 output_declaration_instance322();
    output_declaration323 output_declaration_instance323();
    output_declaration324 output_declaration_instance324();
    output_declaration325 output_declaration_instance325();
    output_declaration326 output_declaration_instance326();
    output_declaration327 output_declaration_instance327();
    output_declaration328 output_declaration_instance328();
    output_declaration329 output_declaration_instance329();
    output_declaration330 output_declaration_instance330();
    output_declaration331 output_declaration_instance331();
    output_declaration332 output_declaration_instance332();
    output_declaration333 output_declaration_instance333();
    output_declaration334 output_declaration_instance334();
    output_declaration335 output_declaration_instance335();
    output_declaration336 output_declaration_instance336();
    output_declaration337 output_declaration_instance337();
    output_declaration338 output_declaration_instance338();
    output_declaration339 output_declaration_instance339();
    output_declaration340 output_declaration_instance340();
    output_declaration341 output_declaration_instance341();
    output_declaration342 output_declaration_instance342();
    output_declaration343 output_declaration_instance343();
    output_declaration344 output_declaration_instance344();
    output_declaration345 output_declaration_instance345();
    output_declaration346 output_declaration_instance346();
    output_declaration347 output_declaration_instance347();
    output_declaration348 output_declaration_instance348();
    output_declaration349 output_declaration_instance349();
    output_declaration350 output_declaration_instance350();
    output_declaration351 output_declaration_instance351();
    output_declaration352 output_declaration_instance352();
    output_declaration353 output_declaration_instance353();
    output_declaration354 output_declaration_instance354();
    output_declaration355 output_declaration_instance355();
    output_declaration356 output_declaration_instance356();
    output_declaration357 output_declaration_instance357();
    output_declaration358 output_declaration_instance358();
    output_declaration359 output_declaration_instance359();
    output_declaration360 output_declaration_instance360();
    output_declaration361 output_declaration_instance361();
    output_declaration362 output_declaration_instance362();
    output_declaration363 output_declaration_instance363();
    output_declaration364 output_declaration_instance364();
    output_declaration365 output_declaration_instance365();
    output_declaration366 output_declaration_instance366();
    output_declaration367 output_declaration_instance367();
    output_declaration368 output_declaration_instance368();
    output_declaration369 output_declaration_instance369();
    output_declaration370 output_declaration_instance370();
    output_declaration371 output_declaration_instance371();
    output_declaration372 output_declaration_instance372();
    output_declaration373 output_declaration_instance373();
    output_declaration374 output_declaration_instance374();
    output_declaration375 output_declaration_instance375();
    output_declaration376 output_declaration_instance376();
    output_declaration377 output_declaration_instance377();
    output_declaration378 output_declaration_instance378();
    output_declaration379 output_declaration_instance379();
    output_declaration380 output_declaration_instance380();
    output_declaration381 output_declaration_instance381();
    output_declaration382 output_declaration_instance382();
    output_declaration383 output_declaration_instance383();
    output_declaration384 output_declaration_instance384();
    output_declaration385 output_declaration_instance385();
    output_declaration386 output_declaration_instance386();
    output_declaration387 output_declaration_instance387();
    output_declaration388 output_declaration_instance388();
    output_declaration389 output_declaration_instance389();
    output_declaration390 output_declaration_instance390();
    output_declaration391 output_declaration_instance391();
    output_declaration392 output_declaration_instance392();
    output_declaration393 output_declaration_instance393();
    output_declaration394 output_declaration_instance394();
    output_declaration395 output_declaration_instance395();
    output_declaration396 output_declaration_instance396();
    output_declaration397 output_declaration_instance397();
    output_declaration398 output_declaration_instance398();
    output_declaration399 output_declaration_instance399();
    output_declaration400 output_declaration_instance400();
    output_declaration401 output_declaration_instance401();
    output_declaration402 output_declaration_instance402();
    output_declaration403 output_declaration_instance403();
    output_declaration404 output_declaration_instance404();
    output_declaration405 output_declaration_instance405();
    output_declaration406 output_declaration_instance406();
    output_declaration407 output_declaration_instance407();
    output_declaration408 output_declaration_instance408();
    output_declaration409 output_declaration_instance409();
    output_declaration410 output_declaration_instance410();
    output_declaration411 output_declaration_instance411();
    output_declaration412 output_declaration_instance412();
    output_declaration413 output_declaration_instance413();
    output_declaration414 output_declaration_instance414();
    output_declaration415 output_declaration_instance415();
    output_declaration416 output_declaration_instance416();
    output_declaration417 output_declaration_instance417();
    output_declaration418 output_declaration_instance418();
    output_declaration419 output_declaration_instance419();
    output_declaration420 output_declaration_instance420();
    output_declaration421 output_declaration_instance421();
    output_declaration422 output_declaration_instance422();
    output_declaration423 output_declaration_instance423();
    output_declaration424 output_declaration_instance424();
    output_declaration425 output_declaration_instance425();
    output_declaration426 output_declaration_instance426();
    output_declaration427 output_declaration_instance427();
    output_declaration428 output_declaration_instance428();
    output_declaration429 output_declaration_instance429();
    output_declaration430 output_declaration_instance430();
    output_declaration431 output_declaration_instance431();
    output_declaration432 output_declaration_instance432();
    output_declaration433 output_declaration_instance433();
    output_declaration434 output_declaration_instance434();
    output_declaration435 output_declaration_instance435();
    output_declaration436 output_declaration_instance436();
    output_declaration437 output_declaration_instance437();
    output_declaration438 output_declaration_instance438();
    output_declaration439 output_declaration_instance439();
    output_declaration440 output_declaration_instance440();
    output_declaration441 output_declaration_instance441();
    output_declaration442 output_declaration_instance442();
    output_declaration443 output_declaration_instance443();
    output_declaration444 output_declaration_instance444();
    output_declaration445 output_declaration_instance445();
    output_declaration446 output_declaration_instance446();
    output_declaration447 output_declaration_instance447();
    output_declaration448 output_declaration_instance448();
    output_declaration449 output_declaration_instance449();
    output_declaration450 output_declaration_instance450();
    output_declaration451 output_declaration_instance451();
    output_declaration452 output_declaration_instance452();
    output_declaration453 output_declaration_instance453();
    output_declaration454 output_declaration_instance454();
    output_declaration455 output_declaration_instance455();
    output_declaration456 output_declaration_instance456();
    output_declaration457 output_declaration_instance457();
    output_declaration458 output_declaration_instance458();
    output_declaration459 output_declaration_instance459();
    output_declaration460 output_declaration_instance460();
    output_declaration461 output_declaration_instance461();
    output_declaration462 output_declaration_instance462();
    output_declaration463 output_declaration_instance463();
    output_declaration464 output_declaration_instance464();
    output_declaration465 output_declaration_instance465();
    output_declaration466 output_declaration_instance466();
    output_declaration467 output_declaration_instance467();
    output_declaration468 output_declaration_instance468();
    output_declaration469 output_declaration_instance469();
    output_declaration470 output_declaration_instance470();
    output_declaration471 output_declaration_instance471();
    output_declaration472 output_declaration_instance472();
    output_declaration473 output_declaration_instance473();
    output_declaration474 output_declaration_instance474();
    output_declaration475 output_declaration_instance475();
    output_declaration476 output_declaration_instance476();
    output_declaration477 output_declaration_instance477();
    output_declaration478 output_declaration_instance478();
    output_declaration479 output_declaration_instance479();
    output_declaration480 output_declaration_instance480();
    output_declaration481 output_declaration_instance481();
    output_declaration482 output_declaration_instance482();
    output_declaration483 output_declaration_instance483();
    output_declaration484 output_declaration_instance484();
    output_declaration485 output_declaration_instance485();
    output_declaration486 output_declaration_instance486();
    output_declaration487 output_declaration_instance487();
    output_declaration488 output_declaration_instance488();
    output_declaration489 output_declaration_instance489();
    output_declaration490 output_declaration_instance490();
    output_declaration491 output_declaration_instance491();
    output_declaration492 output_declaration_instance492();
    output_declaration493 output_declaration_instance493();
    output_declaration494 output_declaration_instance494();
    output_declaration495 output_declaration_instance495();
    output_declaration496 output_declaration_instance496();
    output_declaration497 output_declaration_instance497();
    output_declaration498 output_declaration_instance498();
    output_declaration499 output_declaration_instance499();
    output_declaration500 output_declaration_instance500();
    output_declaration501 output_declaration_instance501();
    output_declaration502 output_declaration_instance502();
    output_declaration503 output_declaration_instance503();
    output_declaration504 output_declaration_instance504();
    output_declaration505 output_declaration_instance505();
    output_declaration506 output_declaration_instance506();
    output_declaration507 output_declaration_instance507();
    output_declaration508 output_declaration_instance508();
    output_declaration509 output_declaration_instance509();
    output_declaration510 output_declaration_instance510();
    output_declaration511 output_declaration_instance511();
    output_declaration512 output_declaration_instance512();
    output_declaration513 output_declaration_instance513();
    output_declaration514 output_declaration_instance514();
    output_declaration515 output_declaration_instance515();
    output_declaration516 output_declaration_instance516();
    output_declaration517 output_declaration_instance517();
    output_declaration518 output_declaration_instance518();
    output_declaration519 output_declaration_instance519();
    output_declaration520 output_declaration_instance520();
    output_declaration521 output_declaration_instance521();
    output_declaration522 output_declaration_instance522();
    output_declaration523 output_declaration_instance523();
    output_declaration524 output_declaration_instance524();
    output_declaration525 output_declaration_instance525();
    output_declaration526 output_declaration_instance526();
    output_declaration527 output_declaration_instance527();
    output_declaration528 output_declaration_instance528();
    output_declaration529 output_declaration_instance529();
    output_declaration530 output_declaration_instance530();
    output_declaration531 output_declaration_instance531();
    output_declaration532 output_declaration_instance532();
    output_declaration533 output_declaration_instance533();
    output_declaration534 output_declaration_instance534();
    output_declaration535 output_declaration_instance535();
    output_declaration536 output_declaration_instance536();
    output_declaration537 output_declaration_instance537();
    output_declaration538 output_declaration_instance538();
    output_declaration539 output_declaration_instance539();
    output_declaration540 output_declaration_instance540();
    output_declaration541 output_declaration_instance541();
    output_declaration542 output_declaration_instance542();
    output_declaration543 output_declaration_instance543();
    output_declaration544 output_declaration_instance544();
    output_declaration545 output_declaration_instance545();
    output_declaration546 output_declaration_instance546();
    output_declaration547 output_declaration_instance547();
    output_declaration548 output_declaration_instance548();
    output_declaration549 output_declaration_instance549();
    output_declaration550 output_declaration_instance550();
    output_declaration551 output_declaration_instance551();
    output_declaration552 output_declaration_instance552();
    output_declaration553 output_declaration_instance553();
    output_declaration554 output_declaration_instance554();
    output_declaration555 output_declaration_instance555();
    output_declaration556 output_declaration_instance556();
    output_declaration557 output_declaration_instance557();
    output_declaration558 output_declaration_instance558();
    output_declaration559 output_declaration_instance559();
    output_declaration560 output_declaration_instance560();
    output_declaration561 output_declaration_instance561();
    output_declaration562 output_declaration_instance562();
    output_declaration563 output_declaration_instance563();
    output_declaration564 output_declaration_instance564();
    output_declaration565 output_declaration_instance565();
    output_declaration566 output_declaration_instance566();
    output_declaration567 output_declaration_instance567();
    output_declaration568 output_declaration_instance568();
    output_declaration569 output_declaration_instance569();
    output_declaration570 output_declaration_instance570();
    output_declaration571 output_declaration_instance571();
    output_declaration572 output_declaration_instance572();
    output_declaration573 output_declaration_instance573();
    output_declaration574 output_declaration_instance574();
    output_declaration575 output_declaration_instance575();
    output_declaration576 output_declaration_instance576();
    output_declaration577 output_declaration_instance577();
    output_declaration578 output_declaration_instance578();
    output_declaration579 output_declaration_instance579();
    output_declaration580 output_declaration_instance580();
    output_declaration581 output_declaration_instance581();
    output_declaration582 output_declaration_instance582();
    output_declaration583 output_declaration_instance583();
    output_declaration584 output_declaration_instance584();
    output_declaration585 output_declaration_instance585();
    output_declaration586 output_declaration_instance586();
    output_declaration587 output_declaration_instance587();
    output_declaration588 output_declaration_instance588();
    output_declaration589 output_declaration_instance589();
    output_declaration590 output_declaration_instance590();
    output_declaration591 output_declaration_instance591();
    output_declaration592 output_declaration_instance592();
    output_declaration593 output_declaration_instance593();
    output_declaration594 output_declaration_instance594();
    output_declaration595 output_declaration_instance595();
    output_declaration596 output_declaration_instance596();
    output_declaration597 output_declaration_instance597();
    output_declaration598 output_declaration_instance598();
    output_declaration599 output_declaration_instance599();
    output_declaration600 output_declaration_instance600();
    output_declaration601 output_declaration_instance601();
    output_declaration602 output_declaration_instance602();
    output_declaration603 output_declaration_instance603();
    output_declaration604 output_declaration_instance604();
    output_declaration605 output_declaration_instance605();
    output_declaration606 output_declaration_instance606();
    output_declaration607 output_declaration_instance607();
    output_declaration608 output_declaration_instance608();
    output_declaration609 output_declaration_instance609();
    output_declaration610 output_declaration_instance610();
    output_declaration611 output_declaration_instance611();
    output_declaration612 output_declaration_instance612();
    output_declaration613 output_declaration_instance613();
    output_declaration614 output_declaration_instance614();
    output_declaration615 output_declaration_instance615();
    output_declaration616 output_declaration_instance616();
    output_declaration617 output_declaration_instance617();
    output_declaration618 output_declaration_instance618();
    output_declaration619 output_declaration_instance619();
    output_declaration620 output_declaration_instance620();
    output_declaration621 output_declaration_instance621();
    output_declaration622 output_declaration_instance622();
    output_declaration623 output_declaration_instance623();
    output_declaration624 output_declaration_instance624();
    output_declaration625 output_declaration_instance625();
    output_declaration626 output_declaration_instance626();
    output_declaration627 output_declaration_instance627();
    output_declaration628 output_declaration_instance628();
    output_declaration629 output_declaration_instance629();
    output_declaration630 output_declaration_instance630();
    output_declaration631 output_declaration_instance631();
    output_declaration632 output_declaration_instance632();
    output_declaration633 output_declaration_instance633();
    output_declaration634 output_declaration_instance634();
    output_declaration635 output_declaration_instance635();
    output_declaration636 output_declaration_instance636();
    output_declaration637 output_declaration_instance637();
    output_declaration638 output_declaration_instance638();
    output_declaration639 output_declaration_instance639();
    output_declaration640 output_declaration_instance640();
    output_declaration641 output_declaration_instance641();
    output_declaration642 output_declaration_instance642();
    output_declaration643 output_declaration_instance643();
    output_declaration644 output_declaration_instance644();
    output_declaration645 output_declaration_instance645();
    output_declaration646 output_declaration_instance646();
    output_declaration647 output_declaration_instance647();
    output_declaration648 output_declaration_instance648();
    output_declaration649 output_declaration_instance649();
    output_declaration650 output_declaration_instance650();
    output_declaration651 output_declaration_instance651();
    output_declaration652 output_declaration_instance652();
    output_declaration653 output_declaration_instance653();
    output_declaration654 output_declaration_instance654();
    output_declaration655 output_declaration_instance655();
    output_declaration656 output_declaration_instance656();
    output_declaration657 output_declaration_instance657();
    output_declaration658 output_declaration_instance658();
    output_declaration659 output_declaration_instance659();
    output_declaration660 output_declaration_instance660();
    output_declaration661 output_declaration_instance661();
    output_declaration662 output_declaration_instance662();
    output_declaration663 output_declaration_instance663();
    output_declaration664 output_declaration_instance664();
    output_declaration665 output_declaration_instance665();
    output_declaration666 output_declaration_instance666();
    output_declaration667 output_declaration_instance667();
    output_declaration668 output_declaration_instance668();
    output_declaration669 output_declaration_instance669();
    output_declaration670 output_declaration_instance670();
    output_declaration671 output_declaration_instance671();
    output_declaration672 output_declaration_instance672();
    output_declaration673 output_declaration_instance673();
    output_declaration674 output_declaration_instance674();
    output_declaration675 output_declaration_instance675();
    output_declaration676 output_declaration_instance676();
    output_declaration677 output_declaration_instance677();
    output_declaration678 output_declaration_instance678();
    output_declaration679 output_declaration_instance679();
    output_declaration680 output_declaration_instance680();
    output_declaration681 output_declaration_instance681();
    output_declaration682 output_declaration_instance682();
    output_declaration683 output_declaration_instance683();
    output_declaration684 output_declaration_instance684();
    output_declaration685 output_declaration_instance685();
    output_declaration686 output_declaration_instance686();
    output_declaration687 output_declaration_instance687();
    output_declaration688 output_declaration_instance688();
    output_declaration689 output_declaration_instance689();
    output_declaration690 output_declaration_instance690();
    output_declaration691 output_declaration_instance691();
    output_declaration692 output_declaration_instance692();
    output_declaration693 output_declaration_instance693();
    output_declaration694 output_declaration_instance694();
    output_declaration695 output_declaration_instance695();
    output_declaration696 output_declaration_instance696();
    output_declaration697 output_declaration_instance697();
    output_declaration698 output_declaration_instance698();
    output_declaration699 output_declaration_instance699();
    output_declaration700 output_declaration_instance700();
    output_declaration701 output_declaration_instance701();
    output_declaration702 output_declaration_instance702();
    output_declaration703 output_declaration_instance703();
    output_declaration704 output_declaration_instance704();
    output_declaration705 output_declaration_instance705();
    output_declaration706 output_declaration_instance706();
    output_declaration707 output_declaration_instance707();
    output_declaration708 output_declaration_instance708();
    output_declaration709 output_declaration_instance709();
    output_declaration710 output_declaration_instance710();
    output_declaration711 output_declaration_instance711();
    output_declaration712 output_declaration_instance712();
    output_declaration713 output_declaration_instance713();
    output_declaration714 output_declaration_instance714();
    output_declaration715 output_declaration_instance715();
    output_declaration716 output_declaration_instance716();
    output_declaration717 output_declaration_instance717();
    output_declaration718 output_declaration_instance718();
    output_declaration719 output_declaration_instance719();
    output_declaration720 output_declaration_instance720();
    output_declaration721 output_declaration_instance721();
    output_declaration722 output_declaration_instance722();
    output_declaration723 output_declaration_instance723();
    output_declaration724 output_declaration_instance724();
    output_declaration725 output_declaration_instance725();
    output_declaration726 output_declaration_instance726();
    output_declaration727 output_declaration_instance727();
    output_declaration728 output_declaration_instance728();
    output_declaration729 output_declaration_instance729();
    output_declaration730 output_declaration_instance730();
    output_declaration731 output_declaration_instance731();
    output_declaration732 output_declaration_instance732();
    output_declaration733 output_declaration_instance733();
    output_declaration734 output_declaration_instance734();
    output_declaration735 output_declaration_instance735();
    output_declaration736 output_declaration_instance736();
    output_declaration737 output_declaration_instance737();
    output_declaration738 output_declaration_instance738();
    output_declaration739 output_declaration_instance739();
    output_declaration740 output_declaration_instance740();
    output_declaration741 output_declaration_instance741();
    output_declaration742 output_declaration_instance742();
    output_declaration743 output_declaration_instance743();
    output_declaration744 output_declaration_instance744();
    output_declaration745 output_declaration_instance745();
    output_declaration746 output_declaration_instance746();
    output_declaration747 output_declaration_instance747();
    output_declaration748 output_declaration_instance748();
    output_declaration749 output_declaration_instance749();
    output_declaration750 output_declaration_instance750();
    output_declaration751 output_declaration_instance751();
    output_declaration752 output_declaration_instance752();
    output_declaration753 output_declaration_instance753();
    output_declaration754 output_declaration_instance754();
    output_declaration755 output_declaration_instance755();
    output_declaration756 output_declaration_instance756();
    output_declaration757 output_declaration_instance757();
    output_declaration758 output_declaration_instance758();
    output_declaration759 output_declaration_instance759();
    output_declaration760 output_declaration_instance760();
    output_declaration761 output_declaration_instance761();
    output_declaration762 output_declaration_instance762();
    output_declaration763 output_declaration_instance763();
    output_declaration764 output_declaration_instance764();
    output_declaration765 output_declaration_instance765();
    output_declaration766 output_declaration_instance766();
    output_declaration767 output_declaration_instance767();
    output_declaration768 output_declaration_instance768();
    output_declaration769 output_declaration_instance769();
    output_declaration770 output_declaration_instance770();
    output_declaration771 output_declaration_instance771();
    output_declaration772 output_declaration_instance772();
    output_declaration773 output_declaration_instance773();
    output_declaration774 output_declaration_instance774();
    output_declaration775 output_declaration_instance775();
    output_declaration776 output_declaration_instance776();
    output_declaration777 output_declaration_instance777();
    output_declaration778 output_declaration_instance778();
    output_declaration779 output_declaration_instance779();
    output_declaration780 output_declaration_instance780();
    output_declaration781 output_declaration_instance781();
    output_declaration782 output_declaration_instance782();
    output_declaration783 output_declaration_instance783();
    output_declaration784 output_declaration_instance784();
    output_declaration785 output_declaration_instance785();
    output_declaration786 output_declaration_instance786();
    output_declaration787 output_declaration_instance787();
    output_declaration788 output_declaration_instance788();
    output_declaration789 output_declaration_instance789();
    output_declaration790 output_declaration_instance790();
    output_declaration791 output_declaration_instance791();
    output_declaration792 output_declaration_instance792();
    output_declaration793 output_declaration_instance793();
    output_declaration794 output_declaration_instance794();
    output_declaration795 output_declaration_instance795();
    output_declaration796 output_declaration_instance796();
    output_declaration797 output_declaration_instance797();
    output_declaration798 output_declaration_instance798();
    output_declaration799 output_declaration_instance799();
    output_declaration800 output_declaration_instance800();
    output_declaration801 output_declaration_instance801();
    output_declaration802 output_declaration_instance802();
    output_declaration803 output_declaration_instance803();
    output_declaration804 output_declaration_instance804();
    output_declaration805 output_declaration_instance805();
    output_declaration806 output_declaration_instance806();
    output_declaration807 output_declaration_instance807();
    output_declaration808 output_declaration_instance808();
    output_declaration809 output_declaration_instance809();
    output_declaration810 output_declaration_instance810();
    output_declaration811 output_declaration_instance811();
    output_declaration812 output_declaration_instance812();
    output_declaration813 output_declaration_instance813();
    output_declaration814 output_declaration_instance814();
    output_declaration815 output_declaration_instance815();
    output_declaration816 output_declaration_instance816();
    output_declaration817 output_declaration_instance817();
    output_declaration818 output_declaration_instance818();
    output_declaration819 output_declaration_instance819();
    output_declaration820 output_declaration_instance820();
    output_declaration821 output_declaration_instance821();
    output_declaration822 output_declaration_instance822();
    output_declaration823 output_declaration_instance823();
    output_declaration824 output_declaration_instance824();
    output_declaration825 output_declaration_instance825();
    output_declaration826 output_declaration_instance826();
    output_declaration827 output_declaration_instance827();
    output_declaration828 output_declaration_instance828();
    output_declaration829 output_declaration_instance829();
    output_declaration830 output_declaration_instance830();
    output_declaration831 output_declaration_instance831();
    output_declaration832 output_declaration_instance832();
    output_declaration833 output_declaration_instance833();
    output_declaration834 output_declaration_instance834();
    output_declaration835 output_declaration_instance835();
    output_declaration836 output_declaration_instance836();
    output_declaration837 output_declaration_instance837();
    output_declaration838 output_declaration_instance838();
    output_declaration839 output_declaration_instance839();
    output_declaration840 output_declaration_instance840();
    output_declaration841 output_declaration_instance841();
    output_declaration842 output_declaration_instance842();
    output_declaration843 output_declaration_instance843();
    output_declaration844 output_declaration_instance844();
    output_declaration845 output_declaration_instance845();
    output_declaration846 output_declaration_instance846();
    output_declaration847 output_declaration_instance847();
    output_declaration848 output_declaration_instance848();
    output_declaration849 output_declaration_instance849();
    output_declaration850 output_declaration_instance850();
    output_declaration851 output_declaration_instance851();
    output_declaration852 output_declaration_instance852();
    output_declaration853 output_declaration_instance853();
    output_declaration854 output_declaration_instance854();
    output_declaration855 output_declaration_instance855();
    output_declaration856 output_declaration_instance856();
    output_declaration857 output_declaration_instance857();
    output_declaration858 output_declaration_instance858();
    output_declaration859 output_declaration_instance859();
    output_declaration860 output_declaration_instance860();
    output_declaration861 output_declaration_instance861();
    output_declaration862 output_declaration_instance862();
    output_declaration863 output_declaration_instance863();
    output_declaration864 output_declaration_instance864();
    output_declaration865 output_declaration_instance865();
    output_declaration866 output_declaration_instance866();
    output_declaration867 output_declaration_instance867();
    output_declaration868 output_declaration_instance868();
    output_declaration869 output_declaration_instance869();
    output_declaration870 output_declaration_instance870();
    output_declaration871 output_declaration_instance871();
    output_declaration872 output_declaration_instance872();
    output_declaration873 output_declaration_instance873();
    output_declaration874 output_declaration_instance874();
    output_declaration875 output_declaration_instance875();
    output_declaration876 output_declaration_instance876();
    output_declaration877 output_declaration_instance877();
    output_declaration878 output_declaration_instance878();
    output_declaration879 output_declaration_instance879();
    output_declaration880 output_declaration_instance880();
    output_declaration881 output_declaration_instance881();
    output_declaration882 output_declaration_instance882();
    output_declaration883 output_declaration_instance883();
    output_declaration884 output_declaration_instance884();
    output_declaration885 output_declaration_instance885();
    output_declaration886 output_declaration_instance886();
    output_declaration887 output_declaration_instance887();
    output_declaration888 output_declaration_instance888();
    output_declaration889 output_declaration_instance889();
    output_declaration890 output_declaration_instance890();
    output_declaration891 output_declaration_instance891();
    output_declaration892 output_declaration_instance892();
    output_declaration893 output_declaration_instance893();
    output_declaration894 output_declaration_instance894();
    output_declaration895 output_declaration_instance895();
endmodule
//@
//author : andreib
module output_declaration0( abc ); output abc;
endmodule
//author : andreib
module output_declaration1( abc ); output [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration2( abc ); output [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration3( abc ); output [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration4( abc ); output [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration5( abc ); output [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration6( abc ); output [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration7( abc ); output [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration8( abc ); output [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration9( abc ); output [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration10( abc ); output [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration11( abc ); output [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration12( abc ); output [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration13( abc ); output [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration14( abc ); output [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration15( abc ); output [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration16( abc ); output [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration17( abc ); output [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration18( abc ); output [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration19( abc ); output [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration20( abc ); output [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration21( abc ); output [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration22( abc ); output [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration23( abc ); output [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration24( abc ); output [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration25( abc ); output [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration26( abc ); output signed abc;
endmodule
//author : andreib
module output_declaration27( abc ); output signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration28( abc ); output signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration29( abc ); output signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration30( abc ); output signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration31( abc ); output signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration32( abc ); output signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration33( abc ); output signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration34( abc ); output signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration35( abc ); output signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration36( abc ); output signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration37( abc ); output signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration38( abc ); output signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration39( abc ); output signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration40( abc ); output signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration41( abc ); output signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration42( abc ); output signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration43( abc ); output signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration44( abc ); output signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration45( abc ); output signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration46( abc ); output signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration47( abc ); output signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration48( abc ); output signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration49( abc ); output signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration50( abc ); output signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration51( abc ); output signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration52( abc ); output supply0 abc;
endmodule
//author : andreib
module output_declaration53( abc ); output supply0 [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration54( abc ); output supply0 [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration55( abc ); output supply0 [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration56( abc ); output supply0 [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration57( abc ); output supply0 [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration58( abc ); output supply0 [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration59( abc ); output supply0 [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration60( abc ); output supply0 [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration61( abc ); output supply0 [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration62( abc ); output supply0 [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration63( abc ); output supply0 [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration64( abc ); output supply0 [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration65( abc ); output supply0 [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration66( abc ); output supply0 [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration67( abc ); output supply0 [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration68( abc ); output supply0 [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration69( abc ); output supply0 [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration70( abc ); output supply0 [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration71( abc ); output supply0 [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration72( abc ); output supply0 [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration73( abc ); output supply0 [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration74( abc ); output supply0 [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration75( abc ); output supply0 [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration76( abc ); output supply0 [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration77( abc ); output supply0 [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration78( abc ); output supply0 signed abc;
endmodule
//author : andreib
module output_declaration79( abc ); output supply0 signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration80( abc ); output supply0 signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration81( abc ); output supply0 signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration82( abc ); output supply0 signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration83( abc ); output supply0 signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration84( abc ); output supply0 signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration85( abc ); output supply0 signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration86( abc ); output supply0 signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration87( abc ); output supply0 signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration88( abc ); output supply0 signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration89( abc ); output supply0 signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration90( abc ); output supply0 signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration91( abc ); output supply0 signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration92( abc ); output supply0 signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration93( abc ); output supply0 signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration94( abc ); output supply0 signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration95( abc ); output supply0 signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration96( abc ); output supply0 signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration97( abc ); output supply0 signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration98( abc ); output supply0 signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration99( abc ); output supply0 signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration100( abc ); output supply0 signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration101( abc ); output supply0 signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration102( abc ); output supply0 signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration103( abc ); output supply0 signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration104( abc ); output supply1 abc;
endmodule
//author : andreib
module output_declaration105( abc ); output supply1 [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration106( abc ); output supply1 [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration107( abc ); output supply1 [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration108( abc ); output supply1 [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration109( abc ); output supply1 [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration110( abc ); output supply1 [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration111( abc ); output supply1 [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration112( abc ); output supply1 [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration113( abc ); output supply1 [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration114( abc ); output supply1 [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration115( abc ); output supply1 [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration116( abc ); output supply1 [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration117( abc ); output supply1 [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration118( abc ); output supply1 [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration119( abc ); output supply1 [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration120( abc ); output supply1 [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration121( abc ); output supply1 [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration122( abc ); output supply1 [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration123( abc ); output supply1 [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration124( abc ); output supply1 [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration125( abc ); output supply1 [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration126( abc ); output supply1 [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration127( abc ); output supply1 [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration128( abc ); output supply1 [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration129( abc ); output supply1 [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration130( abc ); output supply1 signed abc;
endmodule
//author : andreib
module output_declaration131( abc ); output supply1 signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration132( abc ); output supply1 signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration133( abc ); output supply1 signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration134( abc ); output supply1 signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration135( abc ); output supply1 signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration136( abc ); output supply1 signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration137( abc ); output supply1 signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration138( abc ); output supply1 signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration139( abc ); output supply1 signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration140( abc ); output supply1 signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration141( abc ); output supply1 signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration142( abc ); output supply1 signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration143( abc ); output supply1 signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration144( abc ); output supply1 signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration145( abc ); output supply1 signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration146( abc ); output supply1 signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration147( abc ); output supply1 signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration148( abc ); output supply1 signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration149( abc ); output supply1 signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration150( abc ); output supply1 signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration151( abc ); output supply1 signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration152( abc ); output supply1 signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration153( abc ); output supply1 signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration154( abc ); output supply1 signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration155( abc ); output supply1 signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration156( abc ); output tri abc;
endmodule
//author : andreib
module output_declaration157( abc ); output tri [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration158( abc ); output tri [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration159( abc ); output tri [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration160( abc ); output tri [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration161( abc ); output tri [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration162( abc ); output tri [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration163( abc ); output tri [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration164( abc ); output tri [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration165( abc ); output tri [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration166( abc ); output tri [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration167( abc ); output tri [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration168( abc ); output tri [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration169( abc ); output tri [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration170( abc ); output tri [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration171( abc ); output tri [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration172( abc ); output tri [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration173( abc ); output tri [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration174( abc ); output tri [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration175( abc ); output tri [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration176( abc ); output tri [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration177( abc ); output tri [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration178( abc ); output tri [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration179( abc ); output tri [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration180( abc ); output tri [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration181( abc ); output tri [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration182( abc ); output tri signed abc;
endmodule
//author : andreib
module output_declaration183( abc ); output tri signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration184( abc ); output tri signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration185( abc ); output tri signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration186( abc ); output tri signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration187( abc ); output tri signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration188( abc ); output tri signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration189( abc ); output tri signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration190( abc ); output tri signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration191( abc ); output tri signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration192( abc ); output tri signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration193( abc ); output tri signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration194( abc ); output tri signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration195( abc ); output tri signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration196( abc ); output tri signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration197( abc ); output tri signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration198( abc ); output tri signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration199( abc ); output tri signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration200( abc ); output tri signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration201( abc ); output tri signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration202( abc ); output tri signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration203( abc ); output tri signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration204( abc ); output tri signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration205( abc ); output tri signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration206( abc ); output tri signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration207( abc ); output tri signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration208( abc ); output triand abc;
endmodule
//author : andreib
module output_declaration209( abc ); output triand [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration210( abc ); output triand [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration211( abc ); output triand [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration212( abc ); output triand [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration213( abc ); output triand [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration214( abc ); output triand [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration215( abc ); output triand [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration216( abc ); output triand [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration217( abc ); output triand [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration218( abc ); output triand [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration219( abc ); output triand [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration220( abc ); output triand [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration221( abc ); output triand [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration222( abc ); output triand [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration223( abc ); output triand [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration224( abc ); output triand [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration225( abc ); output triand [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration226( abc ); output triand [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration227( abc ); output triand [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration228( abc ); output triand [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration229( abc ); output triand [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration230( abc ); output triand [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration231( abc ); output triand [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration232( abc ); output triand [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration233( abc ); output triand [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration234( abc ); output triand signed abc;
endmodule
//author : andreib
module output_declaration235( abc ); output triand signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration236( abc ); output triand signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration237( abc ); output triand signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration238( abc ); output triand signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration239( abc ); output triand signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration240( abc ); output triand signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration241( abc ); output triand signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration242( abc ); output triand signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration243( abc ); output triand signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration244( abc ); output triand signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration245( abc ); output triand signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration246( abc ); output triand signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration247( abc ); output triand signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration248( abc ); output triand signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration249( abc ); output triand signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration250( abc ); output triand signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration251( abc ); output triand signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration252( abc ); output triand signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration253( abc ); output triand signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration254( abc ); output triand signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration255( abc ); output triand signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration256( abc ); output triand signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration257( abc ); output triand signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration258( abc ); output triand signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration259( abc ); output triand signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration260( abc ); output trior abc;
endmodule
//author : andreib
module output_declaration261( abc ); output trior [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration262( abc ); output trior [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration263( abc ); output trior [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration264( abc ); output trior [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration265( abc ); output trior [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration266( abc ); output trior [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration267( abc ); output trior [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration268( abc ); output trior [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration269( abc ); output trior [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration270( abc ); output trior [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration271( abc ); output trior [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration272( abc ); output trior [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration273( abc ); output trior [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration274( abc ); output trior [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration275( abc ); output trior [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration276( abc ); output trior [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration277( abc ); output trior [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration278( abc ); output trior [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration279( abc ); output trior [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration280( abc ); output trior [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration281( abc ); output trior [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration282( abc ); output trior [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration283( abc ); output trior [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration284( abc ); output trior [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration285( abc ); output trior [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration286( abc ); output trior signed abc;
endmodule
//author : andreib
module output_declaration287( abc ); output trior signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration288( abc ); output trior signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration289( abc ); output trior signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration290( abc ); output trior signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration291( abc ); output trior signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration292( abc ); output trior signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration293( abc ); output trior signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration294( abc ); output trior signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration295( abc ); output trior signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration296( abc ); output trior signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration297( abc ); output trior signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration298( abc ); output trior signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration299( abc ); output trior signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration300( abc ); output trior signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration301( abc ); output trior signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration302( abc ); output trior signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration303( abc ); output trior signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration304( abc ); output trior signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration305( abc ); output trior signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration306( abc ); output trior signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration307( abc ); output trior signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration308( abc ); output trior signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration309( abc ); output trior signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration310( abc ); output trior signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration311( abc ); output trior signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration312( abc ); output tri0 abc;
endmodule
//author : andreib
module output_declaration313( abc ); output tri0 [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration314( abc ); output tri0 [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration315( abc ); output tri0 [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration316( abc ); output tri0 [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration317( abc ); output tri0 [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration318( abc ); output tri0 [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration319( abc ); output tri0 [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration320( abc ); output tri0 [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration321( abc ); output tri0 [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration322( abc ); output tri0 [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration323( abc ); output tri0 [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration324( abc ); output tri0 [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration325( abc ); output tri0 [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration326( abc ); output tri0 [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration327( abc ); output tri0 [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration328( abc ); output tri0 [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration329( abc ); output tri0 [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration330( abc ); output tri0 [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration331( abc ); output tri0 [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration332( abc ); output tri0 [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration333( abc ); output tri0 [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration334( abc ); output tri0 [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration335( abc ); output tri0 [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration336( abc ); output tri0 [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration337( abc ); output tri0 [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration338( abc ); output tri0 signed abc;
endmodule
//author : andreib
module output_declaration339( abc ); output tri0 signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration340( abc ); output tri0 signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration341( abc ); output tri0 signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration342( abc ); output tri0 signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration343( abc ); output tri0 signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration344( abc ); output tri0 signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration345( abc ); output tri0 signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration346( abc ); output tri0 signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration347( abc ); output tri0 signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration348( abc ); output tri0 signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration349( abc ); output tri0 signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration350( abc ); output tri0 signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration351( abc ); output tri0 signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration352( abc ); output tri0 signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration353( abc ); output tri0 signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration354( abc ); output tri0 signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration355( abc ); output tri0 signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration356( abc ); output tri0 signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration357( abc ); output tri0 signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration358( abc ); output tri0 signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration359( abc ); output tri0 signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration360( abc ); output tri0 signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration361( abc ); output tri0 signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration362( abc ); output tri0 signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration363( abc ); output tri0 signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration364( abc ); output tri1 abc;
endmodule
//author : andreib
module output_declaration365( abc ); output tri1 [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration366( abc ); output tri1 [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration367( abc ); output tri1 [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration368( abc ); output tri1 [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration369( abc ); output tri1 [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration370( abc ); output tri1 [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration371( abc ); output tri1 [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration372( abc ); output tri1 [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration373( abc ); output tri1 [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration374( abc ); output tri1 [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration375( abc ); output tri1 [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration376( abc ); output tri1 [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration377( abc ); output tri1 [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration378( abc ); output tri1 [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration379( abc ); output tri1 [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration380( abc ); output tri1 [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration381( abc ); output tri1 [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration382( abc ); output tri1 [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration383( abc ); output tri1 [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration384( abc ); output tri1 [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration385( abc ); output tri1 [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration386( abc ); output tri1 [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration387( abc ); output tri1 [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration388( abc ); output tri1 [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration389( abc ); output tri1 [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration390( abc ); output tri1 signed abc;
endmodule
//author : andreib
module output_declaration391( abc ); output tri1 signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration392( abc ); output tri1 signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration393( abc ); output tri1 signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration394( abc ); output tri1 signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration395( abc ); output tri1 signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration396( abc ); output tri1 signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration397( abc ); output tri1 signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration398( abc ); output tri1 signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration399( abc ); output tri1 signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration400( abc ); output tri1 signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration401( abc ); output tri1 signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration402( abc ); output tri1 signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration403( abc ); output tri1 signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration404( abc ); output tri1 signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration405( abc ); output tri1 signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration406( abc ); output tri1 signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration407( abc ); output tri1 signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration408( abc ); output tri1 signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration409( abc ); output tri1 signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration410( abc ); output tri1 signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration411( abc ); output tri1 signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration412( abc ); output tri1 signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration413( abc ); output tri1 signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration414( abc ); output tri1 signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration415( abc ); output tri1 signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration416( abc ); output wire abc;
endmodule
//author : andreib
module output_declaration417( abc ); output wire [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration418( abc ); output wire [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration419( abc ); output wire [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration420( abc ); output wire [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration421( abc ); output wire [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration422( abc ); output wire [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration423( abc ); output wire [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration424( abc ); output wire [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration425( abc ); output wire [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration426( abc ); output wire [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration427( abc ); output wire [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration428( abc ); output wire [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration429( abc ); output wire [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration430( abc ); output wire [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration431( abc ); output wire [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration432( abc ); output wire [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration433( abc ); output wire [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration434( abc ); output wire [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration435( abc ); output wire [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration436( abc ); output wire [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration437( abc ); output wire [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration438( abc ); output wire [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration439( abc ); output wire [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration440( abc ); output wire [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration441( abc ); output wire [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration442( abc ); output wire signed abc;
endmodule
//author : andreib
module output_declaration443( abc ); output wire signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration444( abc ); output wire signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration445( abc ); output wire signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration446( abc ); output wire signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration447( abc ); output wire signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration448( abc ); output wire signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration449( abc ); output wire signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration450( abc ); output wire signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration451( abc ); output wire signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration452( abc ); output wire signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration453( abc ); output wire signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration454( abc ); output wire signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration455( abc ); output wire signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration456( abc ); output wire signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration457( abc ); output wire signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration458( abc ); output wire signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration459( abc ); output wire signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration460( abc ); output wire signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration461( abc ); output wire signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration462( abc ); output wire signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration463( abc ); output wire signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration464( abc ); output wire signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration465( abc ); output wire signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration466( abc ); output wire signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration467( abc ); output wire signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration468( abc ); output wand abc;
endmodule
//author : andreib
module output_declaration469( abc ); output wand [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration470( abc ); output wand [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration471( abc ); output wand [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration472( abc ); output wand [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration473( abc ); output wand [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration474( abc ); output wand [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration475( abc ); output wand [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration476( abc ); output wand [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration477( abc ); output wand [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration478( abc ); output wand [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration479( abc ); output wand [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration480( abc ); output wand [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration481( abc ); output wand [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration482( abc ); output wand [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration483( abc ); output wand [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration484( abc ); output wand [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration485( abc ); output wand [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration486( abc ); output wand [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration487( abc ); output wand [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration488( abc ); output wand [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration489( abc ); output wand [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration490( abc ); output wand [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration491( abc ); output wand [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration492( abc ); output wand [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration493( abc ); output wand [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration494( abc ); output wand signed abc;
endmodule
//author : andreib
module output_declaration495( abc ); output wand signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration496( abc ); output wand signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration497( abc ); output wand signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration498( abc ); output wand signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration499( abc ); output wand signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration500( abc ); output wand signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration501( abc ); output wand signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration502( abc ); output wand signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration503( abc ); output wand signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration504( abc ); output wand signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration505( abc ); output wand signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration506( abc ); output wand signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration507( abc ); output wand signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration508( abc ); output wand signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration509( abc ); output wand signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration510( abc ); output wand signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration511( abc ); output wand signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration512( abc ); output wand signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration513( abc ); output wand signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration514( abc ); output wand signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration515( abc ); output wand signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration516( abc ); output wand signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration517( abc ); output wand signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration518( abc ); output wand signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration519( abc ); output wand signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration520( abc ); output wor abc;
endmodule
//author : andreib
module output_declaration521( abc ); output wor [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration522( abc ); output wor [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration523( abc ); output wor [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration524( abc ); output wor [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration525( abc ); output wor [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration526( abc ); output wor [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration527( abc ); output wor [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration528( abc ); output wor [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration529( abc ); output wor [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration530( abc ); output wor [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration531( abc ); output wor [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration532( abc ); output wor [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration533( abc ); output wor [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration534( abc ); output wor [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration535( abc ); output wor [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration536( abc ); output wor [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration537( abc ); output wor [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration538( abc ); output wor [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration539( abc ); output wor [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration540( abc ); output wor [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration541( abc ); output wor [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration542( abc ); output wor [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration543( abc ); output wor [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration544( abc ); output wor [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration545( abc ); output wor [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration546( abc ); output wor signed abc;
endmodule
//author : andreib
module output_declaration547( abc ); output wor signed [ 2 : 1 ] abc;
endmodule
//author : andreib
module output_declaration548( abc ); output wor signed [ 2 : +1 ] abc;
endmodule
//author : andreib
module output_declaration549( abc ); output wor signed [ 2 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration550( abc ); output wor signed [ 2 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration551( abc ); output wor signed [ 2 : "str" ] abc;
endmodule
//author : andreib
module output_declaration552( abc ); output wor signed [ +3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration553( abc ); output wor signed [ +3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration554( abc ); output wor signed [ +3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration555( abc ); output wor signed [ +3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration556( abc ); output wor signed [ +3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration557( abc ); output wor signed [ 2-1 : 1 ] abc;
endmodule
//author : andreib
module output_declaration558( abc ); output wor signed [ 2-1 : +1 ] abc;
endmodule
//author : andreib
module output_declaration559( abc ); output wor signed [ 2-1 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration560( abc ); output wor signed [ 2-1 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration561( abc ); output wor signed [ 2-1 : "str" ] abc;
endmodule
//author : andreib
module output_declaration562( abc ); output wor signed [ 1?2:3 : 1 ] abc;
endmodule
//author : andreib
module output_declaration563( abc ); output wor signed [ 1?2:3 : +1 ] abc;
endmodule
//author : andreib
module output_declaration564( abc ); output wor signed [ 1?2:3 : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration565( abc ); output wor signed [ 1?2:3 : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration566( abc ); output wor signed [ 1?2:3 : "str" ] abc;
endmodule
//author : andreib
module output_declaration567( abc ); output wor signed [ "str" : 1 ] abc;
endmodule
//author : andreib
module output_declaration568( abc ); output wor signed [ "str" : +1 ] abc;
endmodule
//author : andreib
module output_declaration569( abc ); output wor signed [ "str" : 2-1 ] abc;
endmodule
//author : andreib
module output_declaration570( abc ); output wor signed [ "str" : 1?2:3 ] abc;
endmodule
//author : andreib
module output_declaration571( abc ); output wor signed [ "str" : "str" ] abc;
endmodule
//author : andreib
module output_declaration572( xyz ); output reg xyz;
endmodule
//author : andreib
module output_declaration573( xyz ); output reg xyz = 2;
endmodule
//author : andreib
module output_declaration574( xyz ); output reg xyz = +3;
endmodule
//author : andreib
module output_declaration575( xyz ); output reg xyz = 2-1;
endmodule
//author : andreib
module output_declaration576( xyz ); output reg xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration577( xyz ); output reg xyz = "str";
endmodule
//author : andreib
module output_declaration578( xyz ); output reg [ 2 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration579( xyz ); output reg [ 2 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration580( xyz ); output reg [ 2 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration581( xyz ); output reg [ 2 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration582( xyz ); output reg [ 2 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration583( xyz ); output reg [ 2 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration584( xyz ); output reg [ 2 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration585( xyz ); output reg [ 2 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration586( xyz ); output reg [ 2 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration587( xyz ); output reg [ 2 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration588( xyz ); output reg [ 2 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration589( xyz ); output reg [ 2 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration590( xyz ); output reg [ 2 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration591( xyz ); output reg [ 2 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration592( xyz ); output reg [ 2 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration593( xyz ); output reg [ 2 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration594( xyz ); output reg [ 2 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration595( xyz ); output reg [ 2 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration596( xyz ); output reg [ 2 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration597( xyz ); output reg [ 2 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration598( xyz ); output reg [ 2 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration599( xyz ); output reg [ 2 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration600( xyz ); output reg [ 2 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration601( xyz ); output reg [ 2 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration602( xyz ); output reg [ 2 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration603( xyz ); output reg [ 2 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration604( xyz ); output reg [ 2 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration605( xyz ); output reg [ 2 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration606( xyz ); output reg [ 2 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration607( xyz ); output reg [ 2 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration608( xyz ); output reg [ +3 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration609( xyz ); output reg [ +3 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration610( xyz ); output reg [ +3 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration611( xyz ); output reg [ +3 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration612( xyz ); output reg [ +3 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration613( xyz ); output reg [ +3 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration614( xyz ); output reg [ +3 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration615( xyz ); output reg [ +3 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration616( xyz ); output reg [ +3 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration617( xyz ); output reg [ +3 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration618( xyz ); output reg [ +3 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration619( xyz ); output reg [ +3 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration620( xyz ); output reg [ +3 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration621( xyz ); output reg [ +3 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration622( xyz ); output reg [ +3 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration623( xyz ); output reg [ +3 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration624( xyz ); output reg [ +3 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration625( xyz ); output reg [ +3 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration626( xyz ); output reg [ +3 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration627( xyz ); output reg [ +3 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration628( xyz ); output reg [ +3 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration629( xyz ); output reg [ +3 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration630( xyz ); output reg [ +3 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration631( xyz ); output reg [ +3 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration632( xyz ); output reg [ +3 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration633( xyz ); output reg [ +3 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration634( xyz ); output reg [ +3 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration635( xyz ); output reg [ +3 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration636( xyz ); output reg [ +3 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration637( xyz ); output reg [ +3 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration638( xyz ); output reg [ 2-1 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration639( xyz ); output reg [ 2-1 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration640( xyz ); output reg [ 2-1 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration641( xyz ); output reg [ 2-1 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration642( xyz ); output reg [ 2-1 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration643( xyz ); output reg [ 2-1 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration644( xyz ); output reg [ 2-1 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration645( xyz ); output reg [ 2-1 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration646( xyz ); output reg [ 2-1 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration647( xyz ); output reg [ 2-1 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration648( xyz ); output reg [ 2-1 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration649( xyz ); output reg [ 2-1 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration650( xyz ); output reg [ 2-1 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration651( xyz ); output reg [ 2-1 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration652( xyz ); output reg [ 2-1 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration653( xyz ); output reg [ 2-1 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration654( xyz ); output reg [ 2-1 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration655( xyz ); output reg [ 2-1 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration656( xyz ); output reg [ 2-1 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration657( xyz ); output reg [ 2-1 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration658( xyz ); output reg [ 2-1 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration659( xyz ); output reg [ 2-1 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration660( xyz ); output reg [ 2-1 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration661( xyz ); output reg [ 2-1 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration662( xyz ); output reg [ 2-1 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration663( xyz ); output reg [ 2-1 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration664( xyz ); output reg [ 2-1 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration665( xyz ); output reg [ 2-1 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration666( xyz ); output reg [ 2-1 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration667( xyz ); output reg [ 2-1 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration668( xyz ); output reg [ 1?2:3 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration669( xyz ); output reg [ 1?2:3 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration670( xyz ); output reg [ 1?2:3 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration671( xyz ); output reg [ 1?2:3 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration672( xyz ); output reg [ 1?2:3 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration673( xyz ); output reg [ 1?2:3 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration674( xyz ); output reg [ 1?2:3 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration675( xyz ); output reg [ 1?2:3 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration676( xyz ); output reg [ 1?2:3 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration677( xyz ); output reg [ 1?2:3 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration678( xyz ); output reg [ 1?2:3 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration679( xyz ); output reg [ 1?2:3 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration680( xyz ); output reg [ 1?2:3 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration681( xyz ); output reg [ 1?2:3 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration682( xyz ); output reg [ 1?2:3 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration683( xyz ); output reg [ 1?2:3 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration684( xyz ); output reg [ 1?2:3 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration685( xyz ); output reg [ 1?2:3 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration686( xyz ); output reg [ 1?2:3 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration687( xyz ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration688( xyz ); output reg [ 1?2:3 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration689( xyz ); output reg [ 1?2:3 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration690( xyz ); output reg [ 1?2:3 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration691( xyz ); output reg [ 1?2:3 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration692( xyz ); output reg [ 1?2:3 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration693( xyz ); output reg [ 1?2:3 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration694( xyz ); output reg [ 1?2:3 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration695( xyz ); output reg [ 1?2:3 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration696( xyz ); output reg [ 1?2:3 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration697( xyz ); output reg [ 1?2:3 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration698( xyz ); output reg [ "str" : 1 ] xyz;
endmodule
//author : andreib
module output_declaration699( xyz ); output reg [ "str" : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration700( xyz ); output reg [ "str" : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration701( xyz ); output reg [ "str" : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration702( xyz ); output reg [ "str" : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration703( xyz ); output reg [ "str" : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration704( xyz ); output reg [ "str" : +1 ] xyz;
endmodule
//author : andreib
module output_declaration705( xyz ); output reg [ "str" : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration706( xyz ); output reg [ "str" : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration707( xyz ); output reg [ "str" : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration708( xyz ); output reg [ "str" : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration709( xyz ); output reg [ "str" : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration710( xyz ); output reg [ "str" : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration711( xyz ); output reg [ "str" : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration712( xyz ); output reg [ "str" : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration713( xyz ); output reg [ "str" : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration714( xyz ); output reg [ "str" : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration715( xyz ); output reg [ "str" : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration716( xyz ); output reg [ "str" : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration717( xyz ); output reg [ "str" : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration718( xyz ); output reg [ "str" : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration719( xyz ); output reg [ "str" : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration720( xyz ); output reg [ "str" : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration721( xyz ); output reg [ "str" : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration722( xyz ); output reg [ "str" : "str" ] xyz;
endmodule
//author : andreib
module output_declaration723( xyz ); output reg [ "str" : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration724( xyz ); output reg [ "str" : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration725( xyz ); output reg [ "str" : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration726( xyz ); output reg [ "str" : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration727( xyz ); output reg [ "str" : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration728( xyz ); output reg signed xyz;
endmodule
//author : andreib
module output_declaration729( xyz ); output reg signed xyz = 2;
endmodule
//author : andreib
module output_declaration730( xyz ); output reg signed xyz = +3;
endmodule
//author : andreib
module output_declaration731( xyz ); output reg signed xyz = 2-1;
endmodule
//author : andreib
module output_declaration732( xyz ); output reg signed xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration733( xyz ); output reg signed xyz = "str";
endmodule
//author : andreib
module output_declaration734( xyz ); output reg signed [ 2 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration735( xyz ); output reg signed [ 2 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration736( xyz ); output reg signed [ 2 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration737( xyz ); output reg signed [ 2 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration738( xyz ); output reg signed [ 2 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration739( xyz ); output reg signed [ 2 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration740( xyz ); output reg signed [ 2 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration741( xyz ); output reg signed [ 2 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration742( xyz ); output reg signed [ 2 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration743( xyz ); output reg signed [ 2 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration744( xyz ); output reg signed [ 2 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration745( xyz ); output reg signed [ 2 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration746( xyz ); output reg signed [ 2 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration747( xyz ); output reg signed [ 2 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration748( xyz ); output reg signed [ 2 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration749( xyz ); output reg signed [ 2 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration750( xyz ); output reg signed [ 2 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration751( xyz ); output reg signed [ 2 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration752( xyz ); output reg signed [ 2 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration753( xyz ); output reg signed [ 2 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration754( xyz ); output reg signed [ 2 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration755( xyz ); output reg signed [ 2 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration756( xyz ); output reg signed [ 2 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration757( xyz ); output reg signed [ 2 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration758( xyz ); output reg signed [ 2 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration759( xyz ); output reg signed [ 2 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration760( xyz ); output reg signed [ 2 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration761( xyz ); output reg signed [ 2 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration762( xyz ); output reg signed [ 2 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration763( xyz ); output reg signed [ 2 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration764( xyz ); output reg signed [ +3 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration765( xyz ); output reg signed [ +3 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration766( xyz ); output reg signed [ +3 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration767( xyz ); output reg signed [ +3 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration768( xyz ); output reg signed [ +3 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration769( xyz ); output reg signed [ +3 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration770( xyz ); output reg signed [ +3 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration771( xyz ); output reg signed [ +3 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration772( xyz ); output reg signed [ +3 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration773( xyz ); output reg signed [ +3 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration774( xyz ); output reg signed [ +3 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration775( xyz ); output reg signed [ +3 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration776( xyz ); output reg signed [ +3 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration777( xyz ); output reg signed [ +3 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration778( xyz ); output reg signed [ +3 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration779( xyz ); output reg signed [ +3 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration780( xyz ); output reg signed [ +3 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration781( xyz ); output reg signed [ +3 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration782( xyz ); output reg signed [ +3 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration783( xyz ); output reg signed [ +3 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration784( xyz ); output reg signed [ +3 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration785( xyz ); output reg signed [ +3 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration786( xyz ); output reg signed [ +3 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration787( xyz ); output reg signed [ +3 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration788( xyz ); output reg signed [ +3 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration789( xyz ); output reg signed [ +3 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration790( xyz ); output reg signed [ +3 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration791( xyz ); output reg signed [ +3 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration792( xyz ); output reg signed [ +3 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration793( xyz ); output reg signed [ +3 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration794( xyz ); output reg signed [ 2-1 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration795( xyz ); output reg signed [ 2-1 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration796( xyz ); output reg signed [ 2-1 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration797( xyz ); output reg signed [ 2-1 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration798( xyz ); output reg signed [ 2-1 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration799( xyz ); output reg signed [ 2-1 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration800( xyz ); output reg signed [ 2-1 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration801( xyz ); output reg signed [ 2-1 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration802( xyz ); output reg signed [ 2-1 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration803( xyz ); output reg signed [ 2-1 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration804( xyz ); output reg signed [ 2-1 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration805( xyz ); output reg signed [ 2-1 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration806( xyz ); output reg signed [ 2-1 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration807( xyz ); output reg signed [ 2-1 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration808( xyz ); output reg signed [ 2-1 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration809( xyz ); output reg signed [ 2-1 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration810( xyz ); output reg signed [ 2-1 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration811( xyz ); output reg signed [ 2-1 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration812( xyz ); output reg signed [ 2-1 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration813( xyz ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration814( xyz ); output reg signed [ 2-1 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration815( xyz ); output reg signed [ 2-1 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration816( xyz ); output reg signed [ 2-1 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration817( xyz ); output reg signed [ 2-1 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration818( xyz ); output reg signed [ 2-1 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration819( xyz ); output reg signed [ 2-1 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration820( xyz ); output reg signed [ 2-1 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration821( xyz ); output reg signed [ 2-1 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration822( xyz ); output reg signed [ 2-1 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration823( xyz ); output reg signed [ 2-1 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration824( xyz ); output reg signed [ 1?2:3 : 1 ] xyz;
endmodule
//author : andreib
module output_declaration825( xyz ); output reg signed [ 1?2:3 : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration826( xyz ); output reg signed [ 1?2:3 : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration827( xyz ); output reg signed [ 1?2:3 : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration828( xyz ); output reg signed [ 1?2:3 : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration829( xyz ); output reg signed [ 1?2:3 : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration830( xyz ); output reg signed [ 1?2:3 : +1 ] xyz;
endmodule
//author : andreib
module output_declaration831( xyz ); output reg signed [ 1?2:3 : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration832( xyz ); output reg signed [ 1?2:3 : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration833( xyz ); output reg signed [ 1?2:3 : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration834( xyz ); output reg signed [ 1?2:3 : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration835( xyz ); output reg signed [ 1?2:3 : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration836( xyz ); output reg signed [ 1?2:3 : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration837( xyz ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration838( xyz ); output reg signed [ 1?2:3 : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration839( xyz ); output reg signed [ 1?2:3 : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration840( xyz ); output reg signed [ 1?2:3 : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration841( xyz ); output reg signed [ 1?2:3 : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration842( xyz ); output reg signed [ 1?2:3 : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration843( xyz ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration844( xyz ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration845( xyz ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration846( xyz ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration847( xyz ); output reg signed [ 1?2:3 : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration848( xyz ); output reg signed [ 1?2:3 : "str" ] xyz;
endmodule
//author : andreib
module output_declaration849( xyz ); output reg signed [ 1?2:3 : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration850( xyz ); output reg signed [ 1?2:3 : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration851( xyz ); output reg signed [ 1?2:3 : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration852( xyz ); output reg signed [ 1?2:3 : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration853( xyz ); output reg signed [ 1?2:3 : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration854( xyz ); output reg signed [ "str" : 1 ] xyz;
endmodule
//author : andreib
module output_declaration855( xyz ); output reg signed [ "str" : 1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration856( xyz ); output reg signed [ "str" : 1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration857( xyz ); output reg signed [ "str" : 1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration858( xyz ); output reg signed [ "str" : 1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration859( xyz ); output reg signed [ "str" : 1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration860( xyz ); output reg signed [ "str" : +1 ] xyz;
endmodule
//author : andreib
module output_declaration861( xyz ); output reg signed [ "str" : +1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration862( xyz ); output reg signed [ "str" : +1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration863( xyz ); output reg signed [ "str" : +1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration864( xyz ); output reg signed [ "str" : +1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration865( xyz ); output reg signed [ "str" : +1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration866( xyz ); output reg signed [ "str" : 2-1 ] xyz;
endmodule
//author : andreib
module output_declaration867( xyz ); output reg signed [ "str" : 2-1 ] xyz = 2;
endmodule
//author : andreib
module output_declaration868( xyz ); output reg signed [ "str" : 2-1 ] xyz = +3;
endmodule
//author : andreib
module output_declaration869( xyz ); output reg signed [ "str" : 2-1 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration870( xyz ); output reg signed [ "str" : 2-1 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration871( xyz ); output reg signed [ "str" : 2-1 ] xyz = "str";
endmodule
//author : andreib
module output_declaration872( xyz ); output reg signed [ "str" : 1?2:3 ] xyz;
endmodule
//author : andreib
module output_declaration873( xyz ); output reg signed [ "str" : 1?2:3 ] xyz = 2;
endmodule
//author : andreib
module output_declaration874( xyz ); output reg signed [ "str" : 1?2:3 ] xyz = +3;
endmodule
//author : andreib
module output_declaration875( xyz ); output reg signed [ "str" : 1?2:3 ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration876( xyz ); output reg signed [ "str" : 1?2:3 ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration877( xyz ); output reg signed [ "str" : 1?2:3 ] xyz = "str";
endmodule
//author : andreib
module output_declaration878( xyz ); output reg signed [ "str" : "str" ] xyz;
endmodule
//author : andreib
module output_declaration879( xyz ); output reg signed [ "str" : "str" ] xyz = 2;
endmodule
//author : andreib
module output_declaration880( xyz ); output reg signed [ "str" : "str" ] xyz = +3;
endmodule
//author : andreib
module output_declaration881( xyz ); output reg signed [ "str" : "str" ] xyz = 2-1;
endmodule
//author : andreib
module output_declaration882( xyz ); output reg signed [ "str" : "str" ] xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration883( xyz ); output reg signed [ "str" : "str" ] xyz = "str";
endmodule
//author : andreib
module output_declaration884( xyz ); output integer xyz;
endmodule
//author : andreib
module output_declaration885( xyz ); output integer xyz = 2;
endmodule
//author : andreib
module output_declaration886( xyz ); output integer xyz = +3;
endmodule
//author : andreib
module output_declaration887( xyz ); output integer xyz = 2-1;
endmodule
//author : andreib
module output_declaration888( xyz ); output integer xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration889( xyz ); output integer xyz = "str";
endmodule
//author : andreib
module output_declaration890( xyz ); output time xyz;
endmodule
//author : andreib
module output_declaration891( xyz ); output time xyz = 2;
endmodule
//author : andreib
module output_declaration892( xyz ); output time xyz = +3;
endmodule
//author : andreib
module output_declaration893( xyz ); output time xyz = 2-1;
endmodule
//author : andreib
module output_declaration894( xyz ); output time xyz = 1?2:3;
endmodule
//author : andreib
module output_declaration895( xyz ); output time xyz = "str";
endmodule
