-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_mbist_cslc_generated/code/vhdl/r_pc.vhd
-- FILE GENERATED ON : Tue Feb 17 20:24:21 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \r_pc\ is
  port(\p_clock\ : in csl_bit;
       \p_reset\ : in csl_bit;
       \p_enable\ : in csl_bit;
       \p_br_addr\ : in csl_bit_vector(10#15# downto 10#0#);
       \p_sel\ : in csl_bit;
       \p_addr_out\ : out csl_bit_vector(10#15# downto 10#0#));
begin
end entity;

architecture \r_pc_logic\ of \r_pc\ is
begin
end architecture;

