`include "defines.v"

module q1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 280
  output [1 - 1:0] ar_sa0_s10;
  p1 p10(.ar_sa0_s10(ar_sa0_s10));
  `include "q1.logic.vh"
endmodule

