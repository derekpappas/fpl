// Test type: initial statement - conditional_statement - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon7;
reg [7:0]a,b;
initial if(a)
	b=0;
endmodule
