-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_cslc_generated/code/vhdl/mem.vhd
-- FILE GENERATED ON : Mon Feb 16 21:37:06 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \mem\ is
  generic(\data_w\ : csl_integer := 10#4#;
          \addr_w\ : csl_integer := 10#8#);
begin
end entity;

architecture \mem_logic\ of \mem\ is
begin
end architecture;

