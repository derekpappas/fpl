-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./proc_ring_cslc_generated/code/vhdl/fabric_drop.vhd
-- FILE GENERATED ON : Wed Jul  9 20:26:20 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \fabric_drop\ is
  port(\db_dwdata\ : out csl_bit_vector(31 downto 0);
       \db_dwwr\ : in csl_bit;
       \dreg_dwdata\ : out csl_bit_vector(31 downto 0);
       \dreg_dwwr\ : in csl_bit;
       \maclu_adwaddr\ : out csl_bit_vector(17 downto 0);
       \maclu_adwdata\ : out csl_bit_vector(31 downto 0);
       \maclu_adwwr\ : in csl_bit;
       \qm_adwaddr\ : out csl_bit_vector(17 downto 0);
       \qm_adwdata\ : out csl_bit_vector(31 downto 0);
       \qm_adwwr\ : in csl_bit;
       \adwraddr\ : out csl_bit_vector(17 downto 0);
       \adwrdata\ : out csl_bit_vector(31 downto 0);
       \adwrwr\ : out csl_bit;
       \adwrrd\ : out csl_bit);
begin
end entity;

architecture \fabric_drop_logic\ of \fabric_drop\ is
begin
end architecture;

