// Test type: Continuous assignment - wk0, sup1 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous196;
wire a;
assign (weak0, supply1) a=1'b1;
endmodule
