`include "defines.v"

module xscalecore();
// Location of source csl unit: file name = IPX2400.csl line number = 259
  `include "xscalecore.logic.v"
endmodule

