--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : b0.vhd
--FILE GENERATED ON : Fri Aug 27 02:46:55 2010


library ieee ; 
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all; 
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
 
use work.csl_util_package.all;

entity b0 is 

 port ( -- Location of source csl unit: file name = temp.csl line number = 7

      ar_sa0_s10: in csl_bit_vector (1 - 1 downto 0)
 );
end b0 ; 

 architecture  arch_b0 of b0 is 
   component a0
     port ( 
      sa0 : in   csl_bit_vector(-1468745200 downto 54) 
 );
  end component; 



 begin
  
a0 : a0 port map ( 
                  sa0 =>(ar_sa0_s10)

              );

 end  arch_b0 ; 
