`include "defines.v"

module m0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 87
  input [1 - 1:0] ar_sa0_s10;
  l0 l0(.ar_sa0_s10(ar_sa0_s10));
  `include "m0.logic.vh"
endmodule

