//test type : task_item_declaration ::= input_declaration
//vparser rule name : 
//author : Codrin
//fixed by: Gabrield
module test_0420;
 task add;
  (* cout = 0, cin = 1 *) input a, b;
  ;
 endtask
endmodule
