//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : i2c.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module i2c(lbdummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 34
  input lbdummy3;
  `include "i2c.logic.v"
endmodule

