include inc8.v
module test;//comm
  `include "../legal/t1.v"
//  /* x */ `include "t1.v"     
//`include "inc0.v"
    endmodule        //end comm
