// Test type: case_statement - casez - default:null
// Vparser rule name:
// Author: andreib
module case_statement48;
reg a;
initial casez(a)
	default: ;
	endcase
endmodule
