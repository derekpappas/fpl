//test type : operator_- concatenation
//vparser rule name : 
//author : Bogdan Mereghea
module unary_operator24;
    wire[1:0] a;
    wire b, c;
    assign a = -{b, c};
endmodule
