`include "defines.v"

module f0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 32
  input [1 - 1:0] ar_sa0_s10;
  e0 e0(.ar_sa0_s10(ar_sa0_s10));
  `include "f0.logic.vh"
endmodule

