`include "defines.v"

module mecluster();
// Location of source csl unit: file name = IPX2400.csl line number = 225
  me me0(), 
     me1(), 
     me2(), 
     me3();
  `include "mecluster.logic.v"
endmodule

