// Test type: Hex Numbers - no size upper case base
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a='H1A3F;
endmodule
