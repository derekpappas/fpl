//cmd_fifo.vh