//gate_instantiation = pulldown ...;
//tests by Gabrield
module gate_instantiation_pulldown0;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown2;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown3;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown4;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown5;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown6;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown7;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown8;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown9;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown10;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown11;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown12;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown13;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown14;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown15;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown16;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown17;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown18;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown19;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown20;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown21;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown22;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown23;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown24;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown25;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown26;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown27;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown28;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown29;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown30;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown31;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown32;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown33;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown34;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown35;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown36;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown37;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown38;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown39;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown40;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown41;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown42;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown43;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown44;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown45;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown46;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown47;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown48;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown49;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown50;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown51;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown52;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown53;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown54;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown55;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown56;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown57;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown58;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown59;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown60;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown61;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown62;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown63;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown64;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown65;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown66;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown67;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown68;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown69;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown70;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown71;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown72;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown73;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown74;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown75;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown76;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown77;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown78;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown79;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown80;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown81;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown82;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown83;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown84;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown85;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown86;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown87;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown88;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown89;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown90;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown91;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown92;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown93;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown94;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown95;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown96;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown97;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown98;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown99;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown100;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown101;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown102;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown103;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown104;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown105;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown106;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown107;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown108;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown109;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown110;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown111;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown112;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown113;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown114;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown115;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown116;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown117;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown118;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown119;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown120;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown121;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown122;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown123;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown124;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown125;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown126;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown127;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown128;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown129;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown130;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown131;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown132;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown133;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown134;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown135;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown136;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown137;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown138;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown139;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown140;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown141;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown142;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown143;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown144;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown145;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown146;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown147;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown148;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown149;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown150;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown151;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown152;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown153;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown154;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown155;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown156;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown157;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown158;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown159;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown160;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown161;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown162;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown163;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown164;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown165;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown166;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown167;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown168;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown169;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown170;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown171;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown172;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown173;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown174;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown175;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown176;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown177;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown178;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown179;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown180;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown181;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown182;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown183;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown184;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown185;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown186;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown187;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown188;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown189;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown190;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown191;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown192;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown193;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown194;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown195;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown196;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown197;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown198;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown199;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown200;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown201;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown202;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown203;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown204;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown205;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown206;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown207;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown208;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown209;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown210;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown211;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown212;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown213;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown214;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown215;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown216;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown217;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown218;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown219;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown220;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown221;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown222;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown223;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown224;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown225;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown226;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown227;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown228;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown229;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown230;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown231;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown232;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown233;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown234;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown235;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown236;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown237;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown238;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown239;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown240;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown241;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown242;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown243;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown244;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown245;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown246;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown247;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown248;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown249;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown250;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown251;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown252;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown253;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown254;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown255;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown256;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown257;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown258;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown259;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown260;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown261;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown262;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown263;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown264;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown265;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown266;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown267;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown268;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown269;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown270;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown271;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown272;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown273;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown274;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown275;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown276;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown277;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown278;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown279;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown280;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown281;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown282;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown283;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown284;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown285;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown286;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown287;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown288;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown289;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown290;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown291;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown292;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown293;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown294;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown295;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown296;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown297;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown298;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown299;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown300;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown301;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown302;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown303;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown304;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown305;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown306;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown307;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown308;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown309;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown310;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown311;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown312;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown313;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown314;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown315;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown316;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown317;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown318;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown319;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown320;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown321;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown322;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown323;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown324;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown325;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown326;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown327;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown328;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown329;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown330;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown331;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown332;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown333;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown334;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown335;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown336;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown337;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown338;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown339;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown340;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown341;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown342;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown343;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown344;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown345;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown346;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown347;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown348;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown349;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown350;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown351;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown352;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown353;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown354;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown355;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown356;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown357;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown358;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown359;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown360;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown361;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown362;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown363;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown364;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown365;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown366;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown367;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown368;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown369;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown370;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown371;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown372;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown373;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown374;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown375;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown376;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown377;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown378;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown379;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown380;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown381;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown382;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown383;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown384;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown385;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown386;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown387;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown388;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown389;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown390;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown391;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown392;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown393;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown394;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown395;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown396;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown397;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown398;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown399;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown400;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown401;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown402;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown403;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown404;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown405;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown406;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown407;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown408;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown409;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown410;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown411;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown412;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown413;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown414;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown415;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown416;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown417;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown418;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown419;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown420;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown421;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown422;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown423;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown424;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown425;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown426;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown427;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown428;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown429;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown430;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown431;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown432;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown433;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown434;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown435;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown436;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown437;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown438;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown439;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown440;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown441;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown442;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown443;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown444;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown445;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown446;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown447;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown448;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown449;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown450;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown451;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown452;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown453;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown454;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown455;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown456;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown457;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown458;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown459;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown460;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown461;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown462;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown463;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown464;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown465;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown466;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown467;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown468;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown469;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown470;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown471;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown472;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown473;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown474;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown475;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown476;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown477;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown478;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown479;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown480;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown481;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown482;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown483;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown484;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown485;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown486;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown487;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown488;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown489;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown490;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown491;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown492;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown493;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown494;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown495;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown496;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown497;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown498;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown499;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown500;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown501;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown502;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown503;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown504;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown505;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown506;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown507;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown508;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown509;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown510;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown511;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown512;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown513;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown514;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown515;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown516;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown517;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown518;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown519;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown520;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown521;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown522;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown523;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown524;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown525;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown526;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown527;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown528;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown529;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown530;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown531;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown532;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown533;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown534;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown535;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown536;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown537;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown538;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown539;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown540;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown541;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown542;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown543;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown544;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown545;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown546;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown547;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown548;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown549;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown550;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown551;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown552;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown553;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown554;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown555;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown556;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown557;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown558;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown559;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown560;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown561;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown562;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown563;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown564;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown565;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown566;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown567;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown568;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown569;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown570;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown571;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown572;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown573;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown574;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown575;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown576;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown577;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown578;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown579;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown580;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown581;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown582;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown583;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown584;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown585;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown586;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown587;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown588;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown589;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown590;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown591;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown592;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown593;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown594;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown595;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown596;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown597;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown598;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown599;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown600;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown601;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown602;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown603;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown604;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown605;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown606;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown607;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown608;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown609;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown610;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown611;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown612;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown613;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown614;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown615;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown616;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown617;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown618;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown619;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown620;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown621;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown622;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown623;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown624;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown625;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown626;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown627;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown628;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown629;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown630;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown631;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown632;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown633;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown634;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown635;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown636;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown637;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown638;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown639;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown640;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown641;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown642;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown643;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown644;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown645;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown646;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown647;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown648;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown649;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown650;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown651;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown652;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown653;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown654;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown655;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown656;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown657;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown658;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown659;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown660;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown661;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown662;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown663;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown664;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown665;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown666;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown667;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown668;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown669;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown670;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown671;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown672;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown673;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown674;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown675;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown676;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown677;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown678;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown679;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown680;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown681;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown682;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown683;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown684;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown685;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown686;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown687;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown688;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown689;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown690;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown691;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown692;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown693;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown694;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown695;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown696;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown697;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown698;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown699;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , supply1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown700;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown701;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown702;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown703;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown704;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown705;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown706;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown707;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown708;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown709;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown710;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown711;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown712;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown713;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown714;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown715;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown716;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown717;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown718;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown719;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown720;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown721;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown722;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown723;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown724;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown725;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown726;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown727;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown728;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown729;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown730;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown731;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown732;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown733;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown734;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown735;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown736;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown737;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown738;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown739;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown740;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown741;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown742;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown743;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown744;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown745;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown746;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown747;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown748;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown749;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , strong1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown750;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown751;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown752;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown753;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown754;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown755;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown756;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown757;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown758;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown759;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown760;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown761;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown762;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown763;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown764;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown765;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown766;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown767;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown768;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown769;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown770;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown771;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown772;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown773;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown774;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown775;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown776;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown777;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown778;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown779;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown780;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown781;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown782;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown783;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown784;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown785;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown786;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown787;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown788;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown789;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown790;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown791;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown792;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown793;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown794;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown795;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown796;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown797;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown798;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown799;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , pull1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown800;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown801;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown802;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown803;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown804;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown805;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown806;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown807;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown808;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown809;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown810;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown811;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown812;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown813;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown814;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown815;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown816;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown817;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown818;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown819;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown820;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown821;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown822;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown823;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown824;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown825;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown826;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown827;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown828;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown829;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown830;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown831;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown832;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown833;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown834;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown835;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown836;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown837;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown838;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown839;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown840;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown841;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown842;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown843;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown844;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown845;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown846;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown847;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown848;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown849;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 , weak1 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown850;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown851;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown852;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown853;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown854;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown855;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown856;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown857;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown858;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown859;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown860;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown861;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown862;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown863;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown864;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown865;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown866;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown867;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown868;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown869;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown870;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown871;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown872;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown873;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown874;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown875;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown876;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown877;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown878;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown879;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown880;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown881;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown882;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown883;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown884;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown885;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown886;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown887;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown888;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown889;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown890;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown891;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown892;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown893;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown894;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown895;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown896;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown897;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown898;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown899;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown900;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown901;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown902;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown903;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown904;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown905;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown906;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown907;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown908;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown909;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown910;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown911;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown912;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown913;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown914;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown915;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown916;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown917;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown918;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown919;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown920;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown921;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown922;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown923;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown924;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown925;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown926;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown927;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown928;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown929;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown930;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown931;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown932;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown933;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown934;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown935;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown936;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown937;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown938;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown939;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown940;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown941;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown942;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown943;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown944;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown945;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown946;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown947;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown948;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown949;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown950;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown951;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown952;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown953;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown954;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown955;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown956;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown957;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown958;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown959;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown960;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown961;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown962;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown963;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown964;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown965;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown966;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown967;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown968;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown969;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown970;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown971;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown972;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown973;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown974;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown975;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown976;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown977;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown978;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown979;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown980;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown981;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown982;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown983;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown984;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown985;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown986;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown987;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown988;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown989;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown990;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown991;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown992;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown993;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown994;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown995;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown996;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown997;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown998;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown999;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1000;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1001;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1002;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1003;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1004;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1005;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1006;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1007;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1008;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1009;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1010;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1011;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1012;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1013;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1014;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1015;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1016;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1017;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1018;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1019;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1020;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1021;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1022;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1023;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1024;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1025;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1026;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1027;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1028;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1029;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1030;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1031;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1032;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1033;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1034;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1035;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1036;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1037;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1038;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1039;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1040;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1041;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1042;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1043;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1044;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1045;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1046;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1047;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1048;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1049;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1050;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1051;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1052;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1053;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1054;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1055;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1056;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1057;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1058;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1059;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1060;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1061;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1062;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1063;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1064;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1065;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1066;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1067;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1068;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1069;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1070;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1071;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1072;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1073;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1074;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1075;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1076;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1077;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1078;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1079;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1080;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1081;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1082;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1083;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1084;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1085;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1086;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1087;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1088;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1089;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1090;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1091;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1092;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1093;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1094;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1095;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1096;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1097;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1098;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1099;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1100;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1101;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1102;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1103;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1104;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1105;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1106;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1107;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1108;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1109;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1110;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1111;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1112;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1113;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1114;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1115;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1116;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1117;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1118;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1119;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1120;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1121;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1122;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1123;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1124;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1125;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1126;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1127;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1128;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1129;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1130;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1131;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1132;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1133;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1134;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1135;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1136;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1137;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1138;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1139;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1140;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1141;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1142;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1143;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1144;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1145;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1146;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1147;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1148;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1149;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1150;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1151;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1152;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1153;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1154;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1155;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1156;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1157;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1158;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1159;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1160;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1161;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1162;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1163;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1164;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1165;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1166;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1167;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1168;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1169;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1170;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1171;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1172;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1173;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1174;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1175;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1176;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1177;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1178;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1179;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1180;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1181;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1182;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1183;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1184;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1185;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1186;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1187;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1188;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1189;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1190;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1191;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1192;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1193;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1194;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1195;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1196;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1197;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1198;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1199;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1200;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1201;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1202;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1203;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1204;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1205;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1206;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1207;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1208;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1209;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1210;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1211;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1212;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1213;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1214;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1215;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1216;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1217;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1218;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1219;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1220;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1221;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1222;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1223;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1224;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1225;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1226;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1227;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1228;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1229;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1230;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1231;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1232;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1233;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1234;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1235;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1236;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1237;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1238;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1239;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1240;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1241;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1242;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1243;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1244;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1245;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1246;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1247;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1248;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1249;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1250;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1251;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1252;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1253;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1254;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1255;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1256;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1257;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1258;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1259;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1260;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1261;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1262;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1263;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1264;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1265;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1266;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1267;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1268;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1269;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1270;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1271;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1272;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1273;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1274;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1275;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1276;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1277;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1278;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1279;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1280;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1281;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1282;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1283;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1284;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1285;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1286;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1287;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1288;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1289;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1290;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1291;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1292;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1293;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1294;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1295;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1296;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1297;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1298;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1299;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1300;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1301;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1302;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1303;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1304;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1305;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1306;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1307;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1308;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1309;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1310;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1311;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1312;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1313;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1314;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1315;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1316;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1317;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1318;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1319;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1320;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1321;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1322;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1323;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1324;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1325;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1326;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1327;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1328;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1329;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1330;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1331;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1332;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1333;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1334;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1335;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1336;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1337;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1338;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1339;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1340;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1341;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1342;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1343;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1344;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1345;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1346;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1347;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1348;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1349;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1350;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1351;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1352;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1353;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1354;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1355;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1356;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1357;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1358;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1359;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1360;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1361;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1362;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1363;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1364;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1365;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1366;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1367;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1368;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1369;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1370;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1371;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1372;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1373;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1374;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1375;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1376;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1377;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1378;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1379;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1380;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1381;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1382;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1383;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1384;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1385;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1386;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1387;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1388;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1389;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1390;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1391;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1392;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1393;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1394;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1395;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1396;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1397;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1398;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1399;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1400;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1401;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1402;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1403;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1404;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1405;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1406;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1407;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1408;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1409;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1410;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1411;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1412;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1413;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1414;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1415;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1416;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1417;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1418;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1419;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1420;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1421;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1422;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1423;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1424;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1425;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1426;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1427;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1428;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1429;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1430;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1431;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1432;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1433;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1434;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1435;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1436;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1437;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1438;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1439;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1440;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1441;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1442;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1443;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1444;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1445;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1446;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1447;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1448;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1449;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1450;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1451;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1452;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1453;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1454;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1455;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1456;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1457;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1458;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1459;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1460;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1461;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1462;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1463;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1464;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1465;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1466;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1467;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1468;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1469;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1470;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1471;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1472;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1473;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1474;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1475;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1476;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1477;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1478;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1479;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1480;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1481;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1482;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1483;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1484;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1485;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1486;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1487;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1488;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1489;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1490;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1491;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1492;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1493;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1494;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1495;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1496;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1497;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1498;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1499;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1500;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1501;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1502;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1503;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1504;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1505;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1506;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1507;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1508;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1509;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1510;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1511;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1512;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1513;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1514;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1515;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1516;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1517;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1518;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1519;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1520;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1521;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1522;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1523;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1524;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1525;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1526;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1527;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1528;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1529;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1530;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1531;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1532;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1533;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1534;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1535;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1536;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1537;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1538;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1539;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1540;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1541;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1542;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1543;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1544;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1545;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1546;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1547;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1548;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1549;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1550;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1551;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1552;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1553;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1554;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1555;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1556;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1557;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1558;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1559;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1560;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1561;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1562;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1563;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1564;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1565;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1566;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1567;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1568;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1569;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1570;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1571;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1572;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1573;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1574;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1575;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1576;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1577;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1578;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1579;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1580;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1581;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1582;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1583;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1584;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1585;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1586;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1587;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1588;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1589;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1590;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1591;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1592;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1593;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1594;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1595;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1596;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1597;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1598;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1599;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1600;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1601;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1602;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1603;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1604;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1605;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1606;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1607;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1608;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1609;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1610;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1611;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1612;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1613;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1614;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1615;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1616;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1617;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1618;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1619;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1620;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1621;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1622;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1623;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1624;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1625;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1626;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1627;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1628;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1629;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1630;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1631;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1632;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1633;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1634;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1635;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1636;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1637;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1638;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1639;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1640;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1641;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1642;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1643;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1644;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1645;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1646;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1647;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1648;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1649;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak1 , weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1650;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1651;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1652;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1653;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1654;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1655;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1656;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1657;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1658;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1659;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1660;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1661;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1662;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1663;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1664;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1665;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1666;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1667;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1668;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1669;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1670;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1671;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1672;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1673;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1674;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1675;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1676;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1677;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1678;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1679;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1680;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1681;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1682;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1683;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1684;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1685;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1686;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1687;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1688;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1689;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1690;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1691;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1692;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1693;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1694;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1695;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1696;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1697;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1698;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1699;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( supply0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1700;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1701;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1702;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1703;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1704;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1705;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1706;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1707;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1708;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1709;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1710;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1711;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1712;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1713;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1714;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1715;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1716;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1717;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1718;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1719;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1720;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1721;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1722;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1723;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1724;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1725;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1726;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1727;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1728;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1729;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1730;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1731;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1732;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1733;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1734;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1735;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1736;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1737;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1738;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1739;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1740;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1741;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1742;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1743;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1744;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1745;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1746;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1747;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1748;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1749;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( strong0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1750;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1751;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1752;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1753;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1754;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1755;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1756;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1757;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1758;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1759;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1760;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1761;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1762;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1763;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1764;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1765;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1766;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1767;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1768;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1769;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1770;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1771;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1772;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1773;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1774;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1775;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1776;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1777;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1778;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1779;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1780;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1781;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1782;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1783;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1784;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1785;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1786;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1787;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1788;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1789;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1790;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1791;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1792;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1793;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1794;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1795;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1796;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1797;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1798;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1799;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( pull0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1800;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1801;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1802;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1803;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1804;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1805;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1806;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1807;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1808;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1809;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1810;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1811;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1812;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1813;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1814;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1815;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1816;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1817;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1818;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1819;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1820;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1821;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1822;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1823;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1824;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( output_terminal ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1825;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1826;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1827;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1828;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1829;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1830;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1831;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1832;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1833;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1834;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1835;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1836;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1837;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1838;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1839;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1840;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1841;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1842;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1843;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1844;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( output_terminal ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1845;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1846;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1847;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , ( multi_output_terminal[7:0] ) ;
endmodule
module gate_instantiation_pulldown1848;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( output_terminal ) ;
endmodule
module gate_instantiation_pulldown1849;
  wire output_terminal;
  wire [7:0] multi_output_terminal;
  pulldown ( weak0 ) ( multi_output_terminal[7:0] ) , name2 ( multi_output_terminal[7:0] ) , name3 ( multi_output_terminal[7:0] ) ;
endmodule
