`include "defines.v"

module e1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 207
  output [1 - 1:0] ar_sa0_s10;
  d1 d10(.ar_sa0_s10(ar_sa0_s10));
  `include "e1.logic.vh"
endmodule

