
module eprom ( cs, rd, address_bus, data_bus, eprom_reset );
input  [15:0] address_bus;
output [15:0] data_bus;
input  cs, rd, eprom_reset;
    wire n147, \mem<2><15> , \mem<4><11> , \mem<8><7> , \mem<7><9> , 
        \mem<12><15> , \mem<2><8> , \mem<2><1> , \mem<6><3> , \mem<11><6> , 
        \mem<3><13> , \mem<13><13> , \n55<9><9> , \mem<2><5> , \mem<3><2> , 
        \mem<9><4> , \mem<7><0> , \mem<10><5> , \mem<9><9> , \mem<11><2> , 
        \mem<2><11> , \mem<6><7> , \mem<12><11> , \mem<3><6> , \mem<4><15> , 
        \mem<7><4> , \mem<8><3> , \mem<10><8> , \mem<10><1> , \mem<3><15> , 
        \mem<5><13> , \mem<9><0> , \mem<5><11> , \mem<9><2> , \mem<11><9> , 
        \mem<13><15> , \mem<7><6> , \mem<3><4> , \mem<8><8> , \mem<10><3> , 
        \mem<2><13> , \mem<12><13> , \mem<2><7> , \mem<8><1> , \mem<11><0> , 
        n_11, \mem<3><0> , \mem<6><5> , \mem<7><2> , \mem<10><7> , 
        \mem<3><11> , \mem<6><8> , \mem<5><15> , \mem<13><11> , \mem<9><6> , 
        \mem<2><3> , \mem<6><1> , \mem<11><4> , \mem<3><9> , \mem<8><5> , 
        \mem<4><13> , \mem<7><12> , \mem<12><8> , \mem<0><5> , \mem<4><7> , 
        \mem<9><10> , \mem<13><2> , \mem<10><10> , n_10, \mem<0><10> , 
        \mem<6><14> , \mem<0><1> , \mem<1><6> , \mem<5><4> , \mem<12><1> , 
        \mem<1><12> , \mem<4><3> , \mem<9><14> , \mem<13><6> , \mem<5><9> , 
        \mem<5><0> , \mem<11><12> , \mem<1><2> , \mem<8><12> , \mem<12><5> , 
        \mem<0><14> , \mem<0><8> , \mem<1><0> , \mem<4><8> , \mem<6><12> , 
        \mem<6><10> , \mem<10><14> , \mem<5><2> , \mem<8><10> , \mem<12><7> , 
        \mem<0><12> , \mem<0><3> , \mem<1><10> , \mem<7><14> , \mem<1><9> , 
        \mem<11><10> , \mem<1><4> , \mem<4><1> , \mem<13><4> , \mem<5><6> , 
        \mem<8><14> , \mem<12><3> , \mem<10><12> , \mem<13><9> , \mem<0><7> , 
        \mem<4><5> , \mem<9><12> , \mem<13><0> , \mem<1><14> , \mem<11><14> , 
        n146, \mem<7><10> , n_15, \mem<0><13> , \mem<1><5> , \mem<12><2> , 
        \mem<5><7> , \mem<8><15> , \mem<10><13> , \mem<13><8> , \mem<0><6> , 
        \mem<4><4> , \mem<9><13> , \mem<13><1> , \mem<11><15> , \mem<1><15> , 
        \mem<7><11> , \mem<1><11> , \mem<1><1> , \mem<4><9> , \mem<6><13> , 
        \mem<5><3> , \mem<8><11> , \mem<12><6> , \mem<7><15> , \mem<0><2> , 
        \mem<1><8> , \mem<11><11> , \mem<13><5> , \mem<0><0> , \mem<4><0> , 
        \mem<9><15> , \mem<13><7> , \mem<1><13> , \mem<4><2> , \mem<5><8> , 
        \n68<0> , \mem<0><15> , \mem<1><3> , \mem<5><1> , \mem<8><13> , 
        \mem<11><13> , \mem<6><11> , \mem<12><4> , \mem<0><9> , \mem<10><15> , 
        \mem<12><9> , n145, \mem<4><6> , \mem<7><13> , n_12, \mem<0><4> , 
        \mem<0><11> , \mem<9><11> , \mem<10><11> , \mem<13><3> , \mem<1><7> , 
        \mem<6><15> , \mem<12><0> , \mem<3><10> , \mem<3><1> , \mem<5><5> , 
        \mem<10><6> , \mem<5><14> , \mem<7><3> , \mem<6><9> , \mem<9><7> , 
        \mem<13><10> , n_13, \mem<2><2> , \mem<6><0> , \mem<3><14> , 
        \mem<3><8> , \mem<11><5> , \mem<4><12> , \mem<8><4> , \mem<9><3> , 
        \mem<13><14> , \mem<11><8> , \mem<3><5> , \mem<5><10> , \mem<7><7> , 
        \mem<8><9> , \mem<8><0> , \mem<10><2> , \mem<12><12> , \mem<2><12> , 
        \mem<2><6> , \mem<11><1> , \mem<2><4> , \mem<6><4> , \mem<9><8> , 
        \mem<11><3> , n_14, \mem<6><6> , \mem<12><10> , \mem<2><14> , 
        \mem<2><10> , \mem<4><14> , \mem<8><2> , \mem<10><9> , \mem<3><7> , 
        \mem<7><5> , \mem<5><12> , \mem<9><1> , \mem<10><0> , \mem<4><10> , 
        \mem<7><8> , \mem<8><6> , \mem<12><14> , \mem<2><9> , \mem<2><0> , 
        \mem<6><2> , \mem<3><12> , \mem<11><7> , \mem<9><5> , \mem<13><12> , 
        \mem<3><3> , \mem<10><4> , \mem<7><1> , n1068, n1067, n1066, n1065, 
        n1064, n1063, n1062, n1061, n1060, n1059, n1058, n1057, n1056, n1055, 
        n1054, n1053, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
        n322, n323, n324, n325, n326, n330, n331, n332, n333, n334, n335, n336, 
        n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
        n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
        n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
        n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
        n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
        n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
        n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
        n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
        n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
        n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
        n457, n458, n459, n684, n727, n728, n729, n730, n731, n732, n733, n734, 
        n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
        n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
        n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
        n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
        n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
        n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
        n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
        n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
        n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, 
        n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
        n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, 
        n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, 
        n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, 
        n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, 
        n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
        n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, 
        n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, 
        n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, 
        n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, 
        n976, n977, n978, n979, n981, n982, n983, n984, n986, n987, n988, n989, 
        n991, n992, n993, n994, n996, n997, n998, n999, n1001, n1002, n1003, 
        n1004, n1006, n1007, n1008, n1009, n1011, n1012, n1013, n1014, n1016, 
        n1017, n1018, n1019, n1021, n1022, n1023, n1024, n1026, n1027, n1028, 
        n1029, n1031, n1032, n1033, n1034, n1036, n1037, n1038, n1039, n1041, 
        n1042, n1043, n1044, n1046, n1047, n1048, n1049, n1051, n1052;
    LD_1 \mem_reg<4><0>  ( .Q(\mem<4><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><13>  ( .Q(\mem<9><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><1>  ( .Q(\mem<13><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><12>  ( .Q(\mem<10><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><2>  ( .Q(\mem<0><2> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<1><15>  ( .Q(\mem<1><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><11>  ( .Q(\mem<7><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><8>  ( .Q(\mem<1><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><1>  ( .Q(\mem<1><1> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<8><15>  ( .Q(\mem<8><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><3>  ( .Q(\mem<5><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><14>  ( .Q(\mem<11><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><13>  ( .Q(\mem<0><13> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<12><2>  ( .Q(\mem<12><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><9>  ( .Q(\mem<4><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><8>  ( .Q(\mem<13><8> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<1><11>  ( .Q(\mem<1><11> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<7><15>  ( .Q(\mem<7><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><6>  ( .Q(\mem<0><6> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<4><4>  ( .Q(\mem<4><4> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<13><5>  ( .Q(\mem<13><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><7>  ( .Q(\mem<5><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><13>  ( .Q(\mem<6><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><6>  ( .Q(\mem<12><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><10>  ( .Q(\mem<11><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><5>  ( .Q(\mem<1><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><11>  ( .Q(\mem<8><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><5>  ( .Q(\mem<5><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><4>  ( .Q(\mem<12><4> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<11><12>  ( .Q(\mem<11><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><7>  ( .Q(\mem<1><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><13>  ( .Q(\mem<8><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><15>  ( .Q(\mem<0><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><11>  ( .Q(\mem<6><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><4>  ( .Q(\mem<0><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><14>  ( .Q(\mem<10><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><6>  ( .Q(\mem<4><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><15>  ( .Q(\mem<9><15> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<13><7>  ( .Q(\mem<13><7> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<0><11>  ( .Q(\mem<0><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><13>  ( .Q(\mem<1><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><9>  ( .Q(\mem<0><9> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<6><15>  ( .Q(\mem<6><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><3>  ( .Q(\mem<1><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><1>  ( .Q(\mem<5><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><0>  ( .Q(\mem<12><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><13>  ( .Q(\mem<7><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><2>  ( .Q(\mem<4><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><8>  ( .Q(\mem<5><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><9>  ( .Q(\mem<12><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><11>  ( .Q(\mem<9><11> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<10><10>  ( .Q(\mem<10><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><3>  ( .Q(\mem<13><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><0>  ( .Q(\mem<0><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><4>  ( .Q(\mem<6><4> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<11><5>  ( .Q(\mem<11><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><11>  ( .Q(\mem<13><11> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<2><6>  ( .Q(\mem<2><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><0>  ( .Q(\mem<8><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><12>  ( .Q(\mem<4><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><5>  ( .Q(\mem<3><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><7>  ( .Q(\mem<7><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><9>  ( .Q(\mem<8><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><6>  ( .Q(\mem<10><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><12>  ( .Q(\mem<2><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><10>  ( .Q(\mem<3><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><14>  ( .Q(\mem<5><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><3>  ( .Q(\mem<9><3> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<3><8>  ( .Q(\mem<3><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><2>  ( .Q(\mem<2><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><4>  ( .Q(\mem<8><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><14>  ( .Q(\mem<3><14> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<6><0>  ( .Q(\mem<6><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><1>  ( .Q(\mem<11><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><15>  ( .Q(\mem<13><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><10>  ( .Q(\mem<5><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><7>  ( .Q(\mem<9><7> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<6><9>  ( .Q(\mem<6><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><8>  ( .Q(\mem<11><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><3>  ( .Q(\mem<7><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><2>  ( .Q(\mem<10><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><13>  ( .Q(\mem<12><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><1>  ( .Q(\mem<3><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><1>  ( .Q(\mem<7><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><0>  ( .Q(\mem<10><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><11>  ( .Q(\mem<12><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><3>  ( .Q(\mem<3><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><12>  ( .Q(\mem<5><12> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<9><5>  ( .Q(\mem<9><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><9>  ( .Q(\mem<2><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><0>  ( .Q(\mem<2><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><10>  ( .Q(\mem<2><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><14>  ( .Q(\mem<4><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><2>  ( .Q(\mem<6><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><3>  ( .Q(\mem<11><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><8>  ( .Q(\mem<7><8> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<10><9>  ( .Q(\mem<10><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><6>  ( .Q(\mem<8><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><12>  ( .Q(\mem<3><12> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<9><1>  ( .Q(\mem<9><1> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<3><7>  ( .Q(\mem<3><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><15>  ( .Q(\mem<12><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><5>  ( .Q(\mem<7><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><4>  ( .Q(\mem<10><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><2>  ( .Q(\mem<8><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><14>  ( .Q(\mem<2><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><10>  ( .Q(\mem<4><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><7>  ( .Q(\mem<11><7> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<6><6>  ( .Q(\mem<6><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><4>  ( .Q(\mem<2><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><8>  ( .Q(\mem<9><8> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<13><13>  ( .Q(\mem<13><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><13>  ( .Q(\mem<3><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><0>  ( .Q(\mem<9><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><6>  ( .Q(\mem<3><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><14>  ( .Q(\mem<12><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><4>  ( .Q(\mem<7><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><5>  ( .Q(\mem<10><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><3>  ( .Q(\mem<8><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><15>  ( .Q(\mem<2><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><11>  ( .Q(\mem<4><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><7>  ( .Q(\mem<6><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><6>  ( .Q(\mem<11><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><12>  ( .Q(\mem<13><12> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<2><5>  ( .Q(\mem<2><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><9>  ( .Q(\mem<9><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><2>  ( .Q(\mem<3><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><0>  ( .Q(\mem<7><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><1>  ( .Q(\mem<10><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><10>  ( .Q(\mem<12><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><8>  ( .Q(\mem<2><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><13>  ( .Q(\mem<5><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><4>  ( .Q(\mem<9><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><1>  ( .Q(\mem<2><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><2>  ( .Q(\mem<11><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><3>  ( .Q(\mem<6><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><9>  ( .Q(\mem<7><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><11>  ( .Q(\mem<2><11> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<10><8>  ( .Q(\mem<10><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><15>  ( .Q(\mem<4><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><7>  ( .Q(\mem<8><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><13>  ( .Q(\mem<2><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><9>  ( .Q(\mem<3><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><5>  ( .Q(\mem<8><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><3>  ( .Q(\mem<2><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><1>  ( .Q(\mem<6><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><0>  ( .Q(\mem<11><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><14>  ( .Q(\mem<13><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><15>  ( .Q(\mem<3><15> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<5><11>  ( .Q(\mem<5><11> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<9><6>  ( .Q(\mem<9><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><8>  ( .Q(\mem<6><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><2>  ( .Q(\mem<7><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><3>  ( .Q(\mem<10><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><9>  ( .Q(\mem<11><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><0>  ( .Q(\mem<3><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><12>  ( .Q(\mem<12><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<2><7>  ( .Q(\mem<2><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><5>  ( .Q(\mem<6><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><4>  ( .Q(\mem<11><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><10>  ( .Q(\mem<13><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><1>  ( .Q(\mem<8><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><13>  ( .Q(\mem<4><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<3><4>  ( .Q(\mem<3><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><8>  ( .Q(\mem<8><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><7>  ( .Q(\mem<10><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><6>  ( .Q(\mem<7><6> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<0><10>  ( .Q(\mem<0><10> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<3><11>  ( .Q(\mem<3><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><15>  ( .Q(\mem<5><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><14>  ( .Q(\mem<6><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><2>  ( .Q(\mem<9><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><8>  ( .Q(\mem<0><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><2>  ( .Q(\mem<1><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><0>  ( .Q(\mem<5><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><1>  ( .Q(\mem<12><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><9>  ( .Q(\mem<5><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><12>  ( .Q(\mem<7><12> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<12><8>  ( .Q(\mem<12><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><1>  ( .Q(\mem<0><1> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<4><3>  ( .Q(\mem<4><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><10>  ( .Q(\mem<9><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><2>  ( .Q(\mem<13><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><11>  ( .Q(\mem<10><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><6>  ( .Q(\mem<1><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><4>  ( .Q(\mem<5><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><13>  ( .Q(\mem<11><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><5>  ( .Q(\mem<12><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><12>  ( .Q(\mem<8><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><14>  ( .Q(\mem<0><14> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<6><10>  ( .Q(\mem<6><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><15>  ( .Q(\mem<10><15> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<0><5>  ( .Q(\mem<0><5> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<4><7>  ( .Q(\mem<4><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><14>  ( .Q(\mem<9><14> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<13><6>  ( .Q(\mem<13><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><12>  ( .Q(\mem<1><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><10>  ( .Q(\mem<1><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<7><14>  ( .Q(\mem<7><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><7>  ( .Q(\mem<0><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><5>  ( .Q(\mem<4><5> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><4>  ( .Q(\mem<13><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<6><12>  ( .Q(\mem<6><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><6>  ( .Q(\mem<5><6> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><11>  ( .Q(\mem<11><11> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><10>  ( .Q(\mem<8><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><7>  ( .Q(\mem<12><7> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><4>  ( .Q(\mem<1><4> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><1>  ( .Q(\mem<4><1> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<9><12>  ( .Q(\mem<9><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><0>  ( .Q(\mem<13><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><3>  ( .Q(\mem<0><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<10><13>  ( .Q(\mem<10><13> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><9>  ( .Q(\mem<1><9> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><14>  ( .Q(\mem<1><14> ), .D(1'b1), .G(n684) );
    LD_1 \mem_reg<7><10>  ( .Q(\mem<7><10> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<1><0>  ( .Q(\mem<1><0> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<8><14>  ( .Q(\mem<8><14> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<5><2>  ( .Q(\mem<5><2> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<12><3>  ( .Q(\mem<12><3> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<0><12>  ( .Q(\mem<0><12> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<4><8>  ( .Q(\mem<4><8> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<11><15>  ( .Q(\mem<11><15> ), .D(1'b0), .G(n684) );
    LD_1 \mem_reg<13><9>  ( .Q(\mem<13><9> ), .D(1'b0), .G(n684) );
    IBUF U539 ( .O(n145), .I(cs) );
    IBUF U540 ( .O(n146), .I(rd) );
    IBUF U541 ( .O(n147), .I(address_bus[15]) );
    IBUF U542 ( .O(n_10), .I(address_bus[5]) );
    IBUF U543 ( .O(n_11), .I(address_bus[4]) );
    IBUF U544 ( .O(n_12), .I(address_bus[3]) );
    IBUF U545 ( .O(n_13), .I(address_bus[2]) );
    IBUF U546 ( .O(n_14), .I(address_bus[1]) );
    IBUF U547 ( .O(n_15), .I(address_bus[0]) );
    OBUF_S U548 ( .O(data_bus[15]), .I(n1053) );
    OBUF_S U549 ( .O(data_bus[14]), .I(n1054) );
    OBUF_S U550 ( .O(data_bus[13]), .I(n1055) );
    OBUF_S U551 ( .O(data_bus[12]), .I(n1056) );
    OBUF_S U552 ( .O(data_bus[11]), .I(n1057) );
    OBUF_S U553 ( .O(data_bus[10]), .I(n1058) );
    OBUF_S U554 ( .O(data_bus[9]), .I(n1059) );
    OBUF_S U555 ( .O(data_bus[8]), .I(n1060) );
    OBUF_S U556 ( .O(data_bus[7]), .I(n1061) );
    OBUF_S U557 ( .O(data_bus[6]), .I(n1062) );
    OBUF_S U558 ( .O(data_bus[5]), .I(n1063) );
    OBUF_S U559 ( .O(data_bus[4]), .I(n1064) );
    OBUF_S U560 ( .O(data_bus[3]), .I(n1065) );
    OBUF_S U561 ( .O(data_bus[2]), .I(n1066) );
    OBUF_S U562 ( .O(data_bus[1]), .I(n1067) );
    OBUF_S U563 ( .O(data_bus[0]), .I(n1068) );
    IBUF U564 ( .O(\n55<9><9> ), .I(eprom_reset) );
    INV U565 ( .O(n684), .I(\n55<9><9> ) );
    OR4 U566 ( .O(n393), .I3(n459), .I2(n458), .I1(n457), .I0(n456) );
    OR4 U567 ( .O(n389), .I3(n455), .I2(n454), .I1(n453), .I0(n452) );
    OR4 U568 ( .O(n385), .I3(n451), .I2(n450), .I1(n449), .I0(n448) );
    OR4 U569 ( .O(n381), .I3(n447), .I2(n446), .I1(n445), .I0(n444) );
    OR4 U570 ( .O(n377), .I3(n443), .I2(n442), .I1(n441), .I0(n440) );
    OR4 U571 ( .O(n373), .I3(n439), .I2(n438), .I1(n437), .I0(n436) );
    OR4 U572 ( .O(n369), .I3(n435), .I2(n434), .I1(n433), .I0(n432) );
    OR4 U573 ( .O(n365), .I3(n431), .I2(n430), .I1(n429), .I0(n428) );
    OR4 U574 ( .O(n361), .I3(n427), .I2(n426), .I1(n425), .I0(n424) );
    OR4 U575 ( .O(n357), .I3(n423), .I2(n422), .I1(n421), .I0(n420) );
    OR4 U576 ( .O(n353), .I3(n419), .I2(n418), .I1(n417), .I0(n416) );
    OR4 U577 ( .O(n349), .I3(n415), .I2(n414), .I1(n413), .I0(n412) );
    OR4 U578 ( .O(n345), .I3(n411), .I2(n410), .I1(n409), .I0(n408) );
    OR4 U579 ( .O(n341), .I3(n407), .I2(n406), .I1(n405), .I0(n404) );
    OR4 U580 ( .O(n337), .I3(n403), .I2(n402), .I1(n401), .I0(n400) );
    OR4 U581 ( .O(n333), .I3(n399), .I2(n398), .I1(n397), .I0(n396) );
    NAND2 U582 ( .O(n728), .I1(\mem<7><0> ), .I0(n319) );
    NAND2 U583 ( .O(n727), .I1(\mem<8><0> ), .I0(n321) );
    NAND2 U584 ( .O(n392), .I1(n727), .I0(n728) );
    NAND2 U585 ( .O(n730), .I1(\mem<9><0> ), .I0(n322) );
    NAND2 U586 ( .O(n729), .I1(\mem<12><0> ), .I0(n325) );
    NAND2 U587 ( .O(n391), .I1(n729), .I0(n730) );
    NAND2 U588 ( .O(n732), .I1(\mem<10><0> ), .I0(n323) );
    NAND2 U589 ( .O(n731), .I1(\mem<13><0> ), .I0(n326) );
    NAND2 U590 ( .O(n390), .I1(n731), .I0(n732) );
    NAND2 U591 ( .O(n734), .I1(\mem<0><0> ), .I0(n314) );
    NAND2 U592 ( .O(n733), .I1(\mem<11><0> ), .I0(n324) );
    NAND2 U593 ( .O(n459), .I1(n733), .I0(n734) );
    NAND2 U594 ( .O(n736), .I1(\mem<1><0> ), .I0(n315) );
    NAND2 U595 ( .O(n735), .I1(n395), .I0(\mem<2><0> ) );
    NAND2 U596 ( .O(n458), .I1(n735), .I0(n736) );
    NAND2 U597 ( .O(n738), .I1(\mem<5><0> ), .I0(n317) );
    NAND2 U598 ( .O(n737), .I1(\mem<6><0> ), .I0(n318) );
    NAND2 U599 ( .O(n457), .I1(n737), .I0(n738) );
    NAND2 U600 ( .O(n740), .I1(\mem<4><0> ), .I0(n316) );
    NAND2 U601 ( .O(n739), .I1(n394), .I0(\mem<3><0> ) );
    NAND2 U602 ( .O(n456), .I1(n739), .I0(n740) );
    NAND2 U603 ( .O(n742), .I1(\mem<7><10> ), .I0(n319) );
    NAND2 U604 ( .O(n741), .I1(\mem<8><10> ), .I0(n321) );
    NAND2 U605 ( .O(n388), .I1(n741), .I0(n742) );
    NAND2 U606 ( .O(n744), .I1(\mem<9><10> ), .I0(n322) );
    NAND2 U607 ( .O(n743), .I1(\mem<12><10> ), .I0(n325) );
    NAND2 U608 ( .O(n387), .I1(n743), .I0(n744) );
    NAND2 U609 ( .O(n746), .I1(\mem<10><10> ), .I0(n323) );
    NAND2 U610 ( .O(n745), .I1(\mem<13><10> ), .I0(n326) );
    NAND2 U611 ( .O(n386), .I1(n745), .I0(n746) );
    NAND2 U612 ( .O(n748), .I1(\mem<0><10> ), .I0(n314) );
    NAND2 U613 ( .O(n747), .I1(\mem<11><10> ), .I0(n324) );
    NAND2 U614 ( .O(n455), .I1(n747), .I0(n748) );
    NAND2 U615 ( .O(n750), .I1(\mem<1><10> ), .I0(n315) );
    NAND2 U616 ( .O(n749), .I1(n395), .I0(\mem<2><10> ) );
    NAND2 U617 ( .O(n454), .I1(n749), .I0(n750) );
    NAND2 U618 ( .O(n752), .I1(\mem<5><10> ), .I0(n317) );
    NAND2 U619 ( .O(n751), .I1(\mem<6><10> ), .I0(n318) );
    NAND2 U620 ( .O(n453), .I1(n751), .I0(n752) );
    NAND2 U621 ( .O(n754), .I1(\mem<4><10> ), .I0(n316) );
    NAND2 U622 ( .O(n753), .I1(n394), .I0(\mem<3><10> ) );
    NAND2 U623 ( .O(n452), .I1(n753), .I0(n754) );
    NAND2 U624 ( .O(n756), .I1(\mem<7><11> ), .I0(n319) );
    NAND2 U625 ( .O(n755), .I1(\mem<8><11> ), .I0(n321) );
    NAND2 U626 ( .O(n384), .I1(n755), .I0(n756) );
    NAND2 U627 ( .O(n758), .I1(\mem<9><11> ), .I0(n322) );
    NAND2 U628 ( .O(n757), .I1(\mem<12><11> ), .I0(n325) );
    NAND2 U629 ( .O(n383), .I1(n757), .I0(n758) );
    NAND2 U630 ( .O(n760), .I1(\mem<10><11> ), .I0(n323) );
    NAND2 U631 ( .O(n759), .I1(\mem<13><11> ), .I0(n326) );
    NAND2 U632 ( .O(n382), .I1(n759), .I0(n760) );
    NAND2 U633 ( .O(n762), .I1(\mem<0><11> ), .I0(n314) );
    NAND2 U634 ( .O(n761), .I1(\mem<11><11> ), .I0(n324) );
    NAND2 U635 ( .O(n451), .I1(n761), .I0(n762) );
    NAND2 U636 ( .O(n764), .I1(\mem<1><11> ), .I0(n315) );
    NAND2 U637 ( .O(n763), .I1(n395), .I0(\mem<2><11> ) );
    NAND2 U638 ( .O(n450), .I1(n763), .I0(n764) );
    NAND2 U639 ( .O(n766), .I1(\mem<5><11> ), .I0(n317) );
    NAND2 U640 ( .O(n765), .I1(\mem<6><11> ), .I0(n318) );
    NAND2 U641 ( .O(n449), .I1(n765), .I0(n766) );
    NAND2 U642 ( .O(n768), .I1(\mem<4><11> ), .I0(n316) );
    NAND2 U643 ( .O(n767), .I1(n394), .I0(\mem<3><11> ) );
    NAND2 U644 ( .O(n448), .I1(n767), .I0(n768) );
    NAND2 U645 ( .O(n770), .I1(\mem<7><12> ), .I0(n319) );
    NAND2 U646 ( .O(n769), .I1(\mem<8><12> ), .I0(n321) );
    NAND2 U647 ( .O(n380), .I1(n769), .I0(n770) );
    NAND2 U648 ( .O(n772), .I1(\mem<9><12> ), .I0(n322) );
    NAND2 U649 ( .O(n771), .I1(\mem<12><12> ), .I0(n325) );
    NAND2 U650 ( .O(n379), .I1(n771), .I0(n772) );
    NAND2 U651 ( .O(n774), .I1(\mem<10><12> ), .I0(n323) );
    NAND2 U652 ( .O(n773), .I1(\mem<13><12> ), .I0(n326) );
    NAND2 U653 ( .O(n378), .I1(n773), .I0(n774) );
    NAND2 U654 ( .O(n776), .I1(\mem<0><12> ), .I0(n314) );
    NAND2 U655 ( .O(n775), .I1(\mem<11><12> ), .I0(n324) );
    NAND2 U656 ( .O(n447), .I1(n775), .I0(n776) );
    NAND2 U657 ( .O(n778), .I1(\mem<1><12> ), .I0(n315) );
    NAND2 U658 ( .O(n777), .I1(n395), .I0(\mem<2><12> ) );
    NAND2 U659 ( .O(n446), .I1(n777), .I0(n778) );
    NAND2 U660 ( .O(n780), .I1(\mem<5><12> ), .I0(n317) );
    NAND2 U661 ( .O(n779), .I1(\mem<6><12> ), .I0(n318) );
    NAND2 U662 ( .O(n445), .I1(n779), .I0(n780) );
    NAND2 U663 ( .O(n782), .I1(\mem<4><12> ), .I0(n316) );
    NAND2 U664 ( .O(n781), .I1(n394), .I0(\mem<3><12> ) );
    NAND2 U665 ( .O(n444), .I1(n781), .I0(n782) );
    NAND2 U666 ( .O(n784), .I1(\mem<7><13> ), .I0(n319) );
    NAND2 U667 ( .O(n783), .I1(\mem<8><13> ), .I0(n321) );
    NAND2 U668 ( .O(n376), .I1(n783), .I0(n784) );
    NAND2 U669 ( .O(n786), .I1(\mem<9><13> ), .I0(n322) );
    NAND2 U670 ( .O(n785), .I1(\mem<12><13> ), .I0(n325) );
    NAND2 U671 ( .O(n375), .I1(n785), .I0(n786) );
    NAND2 U672 ( .O(n788), .I1(\mem<10><13> ), .I0(n323) );
    NAND2 U673 ( .O(n787), .I1(\mem<13><13> ), .I0(n326) );
    NAND2 U674 ( .O(n374), .I1(n787), .I0(n788) );
    NAND2 U675 ( .O(n790), .I1(\mem<0><13> ), .I0(n314) );
    NAND2 U676 ( .O(n789), .I1(\mem<11><13> ), .I0(n324) );
    NAND2 U677 ( .O(n443), .I1(n789), .I0(n790) );
    NAND2 U678 ( .O(n792), .I1(\mem<1><13> ), .I0(n315) );
    NAND2 U679 ( .O(n791), .I1(n395), .I0(\mem<2><13> ) );
    NAND2 U680 ( .O(n442), .I1(n791), .I0(n792) );
    NAND2 U681 ( .O(n794), .I1(\mem<5><13> ), .I0(n317) );
    NAND2 U682 ( .O(n793), .I1(\mem<6><13> ), .I0(n318) );
    NAND2 U683 ( .O(n441), .I1(n793), .I0(n794) );
    NAND2 U684 ( .O(n796), .I1(\mem<4><13> ), .I0(n316) );
    NAND2 U685 ( .O(n795), .I1(n394), .I0(\mem<3><13> ) );
    NAND2 U686 ( .O(n440), .I1(n795), .I0(n796) );
    NAND2 U687 ( .O(n798), .I1(\mem<7><14> ), .I0(n319) );
    NAND2 U688 ( .O(n797), .I1(\mem<8><14> ), .I0(n321) );
    NAND2 U689 ( .O(n372), .I1(n797), .I0(n798) );
    NAND2 U690 ( .O(n800), .I1(\mem<9><14> ), .I0(n322) );
    NAND2 U691 ( .O(n799), .I1(\mem<12><14> ), .I0(n325) );
    NAND2 U692 ( .O(n371), .I1(n799), .I0(n800) );
    NAND2 U693 ( .O(n802), .I1(\mem<10><14> ), .I0(n323) );
    NAND2 U694 ( .O(n801), .I1(\mem<13><14> ), .I0(n326) );
    NAND2 U695 ( .O(n370), .I1(n801), .I0(n802) );
    NAND2 U696 ( .O(n804), .I1(\mem<0><14> ), .I0(n314) );
    NAND2 U697 ( .O(n803), .I1(\mem<11><14> ), .I0(n324) );
    NAND2 U698 ( .O(n439), .I1(n803), .I0(n804) );
    NAND2 U699 ( .O(n806), .I1(\mem<1><14> ), .I0(n315) );
    NAND2 U700 ( .O(n805), .I1(n395), .I0(\mem<2><14> ) );
    NAND2 U701 ( .O(n438), .I1(n805), .I0(n806) );
    NAND2 U702 ( .O(n808), .I1(\mem<5><14> ), .I0(n317) );
    NAND2 U703 ( .O(n807), .I1(\mem<6><14> ), .I0(n318) );
    NAND2 U704 ( .O(n437), .I1(n807), .I0(n808) );
    NAND2 U705 ( .O(n810), .I1(\mem<4><14> ), .I0(n316) );
    NAND2 U706 ( .O(n809), .I1(n394), .I0(\mem<3><14> ) );
    NAND2 U707 ( .O(n436), .I1(n809), .I0(n810) );
    NAND2 U708 ( .O(n812), .I1(\mem<7><15> ), .I0(n319) );
    NAND2 U709 ( .O(n811), .I1(\mem<8><15> ), .I0(n321) );
    NAND2 U710 ( .O(n368), .I1(n811), .I0(n812) );
    NAND2 U711 ( .O(n814), .I1(\mem<9><15> ), .I0(n322) );
    NAND2 U712 ( .O(n813), .I1(\mem<12><15> ), .I0(n325) );
    NAND2 U713 ( .O(n367), .I1(n813), .I0(n814) );
    NAND2 U714 ( .O(n816), .I1(\mem<10><15> ), .I0(n323) );
    NAND2 U715 ( .O(n815), .I1(\mem<13><15> ), .I0(n326) );
    NAND2 U716 ( .O(n366), .I1(n815), .I0(n816) );
    NAND2 U717 ( .O(n818), .I1(\mem<0><15> ), .I0(n314) );
    NAND2 U718 ( .O(n817), .I1(\mem<11><15> ), .I0(n324) );
    NAND2 U719 ( .O(n435), .I1(n817), .I0(n818) );
    NAND2 U720 ( .O(n820), .I1(\mem<1><15> ), .I0(n315) );
    NAND2 U721 ( .O(n819), .I1(n395), .I0(\mem<2><15> ) );
    NAND2 U722 ( .O(n434), .I1(n819), .I0(n820) );
    NAND2 U723 ( .O(n822), .I1(\mem<5><15> ), .I0(n317) );
    NAND2 U724 ( .O(n821), .I1(\mem<6><15> ), .I0(n318) );
    NAND2 U725 ( .O(n433), .I1(n821), .I0(n822) );
    NAND2 U726 ( .O(n824), .I1(\mem<4><15> ), .I0(n316) );
    NAND2 U727 ( .O(n823), .I1(n394), .I0(\mem<3><15> ) );
    NAND2 U728 ( .O(n432), .I1(n823), .I0(n824) );
    NAND2 U729 ( .O(n826), .I1(\mem<7><1> ), .I0(n319) );
    NAND2 U730 ( .O(n825), .I1(\mem<8><1> ), .I0(n321) );
    NAND2 U731 ( .O(n364), .I1(n825), .I0(n826) );
    NAND2 U732 ( .O(n828), .I1(\mem<9><1> ), .I0(n322) );
    NAND2 U733 ( .O(n827), .I1(\mem<12><1> ), .I0(n325) );
    NAND2 U734 ( .O(n363), .I1(n827), .I0(n828) );
    NAND2 U735 ( .O(n830), .I1(\mem<10><1> ), .I0(n323) );
    NAND2 U736 ( .O(n829), .I1(\mem<13><1> ), .I0(n326) );
    NAND2 U737 ( .O(n362), .I1(n829), .I0(n830) );
    NAND2 U738 ( .O(n832), .I1(\mem<0><1> ), .I0(n314) );
    NAND2 U739 ( .O(n831), .I1(\mem<11><1> ), .I0(n324) );
    NAND2 U740 ( .O(n431), .I1(n831), .I0(n832) );
    NAND2 U741 ( .O(n834), .I1(\mem<1><1> ), .I0(n315) );
    NAND2 U742 ( .O(n833), .I1(n395), .I0(\mem<2><1> ) );
    NAND2 U743 ( .O(n430), .I1(n833), .I0(n834) );
    NAND2 U744 ( .O(n836), .I1(\mem<5><1> ), .I0(n317) );
    NAND2 U745 ( .O(n835), .I1(\mem<6><1> ), .I0(n318) );
    NAND2 U746 ( .O(n429), .I1(n835), .I0(n836) );
    NAND2 U747 ( .O(n838), .I1(\mem<4><1> ), .I0(n316) );
    NAND2 U748 ( .O(n837), .I1(n394), .I0(\mem<3><1> ) );
    NAND2 U749 ( .O(n428), .I1(n837), .I0(n838) );
    NAND2 U750 ( .O(n840), .I1(\mem<7><2> ), .I0(n319) );
    NAND2 U751 ( .O(n839), .I1(\mem<8><2> ), .I0(n321) );
    NAND2 U752 ( .O(n360), .I1(n839), .I0(n840) );
    NAND2 U753 ( .O(n842), .I1(\mem<9><2> ), .I0(n322) );
    NAND2 U754 ( .O(n841), .I1(\mem<12><2> ), .I0(n325) );
    NAND2 U755 ( .O(n359), .I1(n841), .I0(n842) );
    NAND2 U756 ( .O(n844), .I1(\mem<10><2> ), .I0(n323) );
    NAND2 U757 ( .O(n843), .I1(\mem<13><2> ), .I0(n326) );
    NAND2 U758 ( .O(n358), .I1(n843), .I0(n844) );
    NAND2 U759 ( .O(n846), .I1(\mem<0><2> ), .I0(n314) );
    NAND2 U760 ( .O(n845), .I1(\mem<11><2> ), .I0(n324) );
    NAND2 U761 ( .O(n427), .I1(n845), .I0(n846) );
    NAND2 U762 ( .O(n848), .I1(\mem<1><2> ), .I0(n315) );
    NAND2 U763 ( .O(n847), .I1(n395), .I0(\mem<2><2> ) );
    NAND2 U764 ( .O(n426), .I1(n847), .I0(n848) );
    NAND2 U765 ( .O(n850), .I1(\mem<5><2> ), .I0(n317) );
    NAND2 U766 ( .O(n849), .I1(\mem<6><2> ), .I0(n318) );
    NAND2 U767 ( .O(n425), .I1(n849), .I0(n850) );
    NAND2 U768 ( .O(n852), .I1(\mem<4><2> ), .I0(n316) );
    NAND2 U769 ( .O(n851), .I1(n394), .I0(\mem<3><2> ) );
    NAND2 U770 ( .O(n424), .I1(n851), .I0(n852) );
    NAND2 U771 ( .O(n854), .I1(\mem<7><3> ), .I0(n319) );
    NAND2 U772 ( .O(n853), .I1(\mem<8><3> ), .I0(n321) );
    NAND2 U773 ( .O(n356), .I1(n853), .I0(n854) );
    NAND2 U774 ( .O(n856), .I1(\mem<9><3> ), .I0(n322) );
    NAND2 U775 ( .O(n855), .I1(\mem<12><3> ), .I0(n325) );
    NAND2 U776 ( .O(n355), .I1(n855), .I0(n856) );
    NAND2 U777 ( .O(n858), .I1(\mem<10><3> ), .I0(n323) );
    NAND2 U778 ( .O(n857), .I1(\mem<13><3> ), .I0(n326) );
    NAND2 U779 ( .O(n354), .I1(n857), .I0(n858) );
    NAND2 U780 ( .O(n860), .I1(\mem<0><3> ), .I0(n314) );
    NAND2 U781 ( .O(n859), .I1(\mem<11><3> ), .I0(n324) );
    NAND2 U782 ( .O(n423), .I1(n859), .I0(n860) );
    NAND2 U783 ( .O(n862), .I1(\mem<1><3> ), .I0(n315) );
    NAND2 U784 ( .O(n861), .I1(n395), .I0(\mem<2><3> ) );
    NAND2 U785 ( .O(n422), .I1(n861), .I0(n862) );
    NAND2 U786 ( .O(n864), .I1(\mem<5><3> ), .I0(n317) );
    NAND2 U787 ( .O(n863), .I1(\mem<6><3> ), .I0(n318) );
    NAND2 U788 ( .O(n421), .I1(n863), .I0(n864) );
    NAND2 U789 ( .O(n866), .I1(\mem<4><3> ), .I0(n316) );
    NAND2 U790 ( .O(n865), .I1(n394), .I0(\mem<3><3> ) );
    NAND2 U791 ( .O(n420), .I1(n865), .I0(n866) );
    NAND2 U792 ( .O(n868), .I1(\mem<7><4> ), .I0(n319) );
    NAND2 U793 ( .O(n867), .I1(\mem<8><4> ), .I0(n321) );
    NAND2 U794 ( .O(n352), .I1(n867), .I0(n868) );
    NAND2 U795 ( .O(n870), .I1(\mem<9><4> ), .I0(n322) );
    NAND2 U796 ( .O(n869), .I1(\mem<12><4> ), .I0(n325) );
    NAND2 U797 ( .O(n351), .I1(n869), .I0(n870) );
    NAND2 U798 ( .O(n872), .I1(\mem<10><4> ), .I0(n323) );
    NAND2 U799 ( .O(n871), .I1(\mem<13><4> ), .I0(n326) );
    NAND2 U800 ( .O(n350), .I1(n871), .I0(n872) );
    NAND2 U801 ( .O(n874), .I1(\mem<0><4> ), .I0(n314) );
    NAND2 U802 ( .O(n873), .I1(\mem<11><4> ), .I0(n324) );
    NAND2 U803 ( .O(n419), .I1(n873), .I0(n874) );
    NAND2 U804 ( .O(n876), .I1(\mem<1><4> ), .I0(n315) );
    NAND2 U805 ( .O(n875), .I1(n395), .I0(\mem<2><4> ) );
    NAND2 U806 ( .O(n418), .I1(n875), .I0(n876) );
    NAND2 U807 ( .O(n878), .I1(\mem<5><4> ), .I0(n317) );
    NAND2 U808 ( .O(n877), .I1(\mem<6><4> ), .I0(n318) );
    NAND2 U809 ( .O(n417), .I1(n877), .I0(n878) );
    NAND2 U810 ( .O(n880), .I1(\mem<4><4> ), .I0(n316) );
    NAND2 U811 ( .O(n879), .I1(n394), .I0(\mem<3><4> ) );
    NAND2 U812 ( .O(n416), .I1(n879), .I0(n880) );
    NAND2 U813 ( .O(n882), .I1(\mem<7><5> ), .I0(n319) );
    NAND2 U814 ( .O(n881), .I1(\mem<8><5> ), .I0(n321) );
    NAND2 U815 ( .O(n348), .I1(n881), .I0(n882) );
    NAND2 U816 ( .O(n884), .I1(\mem<9><5> ), .I0(n322) );
    NAND2 U817 ( .O(n883), .I1(\mem<12><5> ), .I0(n325) );
    NAND2 U818 ( .O(n347), .I1(n883), .I0(n884) );
    NAND2 U819 ( .O(n886), .I1(\mem<10><5> ), .I0(n323) );
    NAND2 U820 ( .O(n885), .I1(\mem<13><5> ), .I0(n326) );
    NAND2 U821 ( .O(n346), .I1(n885), .I0(n886) );
    NAND2 U822 ( .O(n888), .I1(\mem<0><5> ), .I0(n314) );
    NAND2 U823 ( .O(n887), .I1(\mem<11><5> ), .I0(n324) );
    NAND2 U824 ( .O(n415), .I1(n887), .I0(n888) );
    NAND2 U825 ( .O(n890), .I1(\mem<1><5> ), .I0(n315) );
    NAND2 U826 ( .O(n889), .I1(n395), .I0(\mem<2><5> ) );
    NAND2 U827 ( .O(n414), .I1(n889), .I0(n890) );
    NAND2 U828 ( .O(n892), .I1(\mem<5><5> ), .I0(n317) );
    NAND2 U829 ( .O(n891), .I1(\mem<6><5> ), .I0(n318) );
    NAND2 U830 ( .O(n413), .I1(n891), .I0(n892) );
    NAND2 U831 ( .O(n894), .I1(\mem<4><5> ), .I0(n316) );
    NAND2 U832 ( .O(n893), .I1(n394), .I0(\mem<3><5> ) );
    NAND2 U833 ( .O(n412), .I1(n893), .I0(n894) );
    NAND2 U834 ( .O(n896), .I1(\mem<7><6> ), .I0(n319) );
    NAND2 U835 ( .O(n895), .I1(\mem<8><6> ), .I0(n321) );
    NAND2 U836 ( .O(n344), .I1(n895), .I0(n896) );
    NAND2 U837 ( .O(n898), .I1(\mem<9><6> ), .I0(n322) );
    NAND2 U838 ( .O(n897), .I1(\mem<12><6> ), .I0(n325) );
    NAND2 U839 ( .O(n343), .I1(n897), .I0(n898) );
    NAND2 U840 ( .O(n900), .I1(\mem<10><6> ), .I0(n323) );
    NAND2 U841 ( .O(n899), .I1(\mem<13><6> ), .I0(n326) );
    NAND2 U842 ( .O(n342), .I1(n899), .I0(n900) );
    NAND2 U843 ( .O(n902), .I1(\mem<0><6> ), .I0(n314) );
    NAND2 U844 ( .O(n901), .I1(\mem<11><6> ), .I0(n324) );
    NAND2 U845 ( .O(n411), .I1(n901), .I0(n902) );
    NAND2 U846 ( .O(n904), .I1(\mem<1><6> ), .I0(n315) );
    NAND2 U847 ( .O(n903), .I1(n395), .I0(\mem<2><6> ) );
    NAND2 U848 ( .O(n410), .I1(n903), .I0(n904) );
    NAND2 U849 ( .O(n906), .I1(\mem<5><6> ), .I0(n317) );
    NAND2 U850 ( .O(n905), .I1(\mem<6><6> ), .I0(n318) );
    NAND2 U851 ( .O(n409), .I1(n905), .I0(n906) );
    NAND2 U852 ( .O(n908), .I1(\mem<4><6> ), .I0(n316) );
    NAND2 U853 ( .O(n907), .I1(n394), .I0(\mem<3><6> ) );
    NAND2 U854 ( .O(n408), .I1(n907), .I0(n908) );
    NAND2 U855 ( .O(n910), .I1(\mem<7><7> ), .I0(n319) );
    NAND2 U856 ( .O(n909), .I1(\mem<8><7> ), .I0(n321) );
    NAND2 U857 ( .O(n340), .I1(n909), .I0(n910) );
    NAND2 U858 ( .O(n912), .I1(\mem<9><7> ), .I0(n322) );
    NAND2 U859 ( .O(n911), .I1(\mem<12><7> ), .I0(n325) );
    NAND2 U860 ( .O(n339), .I1(n911), .I0(n912) );
    NAND2 U861 ( .O(n914), .I1(\mem<10><7> ), .I0(n323) );
    NAND2 U862 ( .O(n913), .I1(\mem<13><7> ), .I0(n326) );
    NAND2 U863 ( .O(n338), .I1(n913), .I0(n914) );
    NAND2 U864 ( .O(n916), .I1(\mem<0><7> ), .I0(n314) );
    NAND2 U865 ( .O(n915), .I1(\mem<11><7> ), .I0(n324) );
    NAND2 U866 ( .O(n407), .I1(n915), .I0(n916) );
    NAND2 U867 ( .O(n918), .I1(\mem<1><7> ), .I0(n315) );
    NAND2 U868 ( .O(n917), .I1(n395), .I0(\mem<2><7> ) );
    NAND2 U869 ( .O(n406), .I1(n917), .I0(n918) );
    NAND2 U870 ( .O(n920), .I1(\mem<5><7> ), .I0(n317) );
    NAND2 U871 ( .O(n919), .I1(\mem<6><7> ), .I0(n318) );
    NAND2 U872 ( .O(n405), .I1(n919), .I0(n920) );
    NAND2 U873 ( .O(n922), .I1(\mem<4><7> ), .I0(n316) );
    NAND2 U874 ( .O(n921), .I1(n394), .I0(\mem<3><7> ) );
    NAND2 U875 ( .O(n404), .I1(n921), .I0(n922) );
    NAND2 U876 ( .O(n924), .I1(\mem<7><8> ), .I0(n319) );
    NAND2 U877 ( .O(n923), .I1(\mem<8><8> ), .I0(n321) );
    NAND2 U878 ( .O(n336), .I1(n923), .I0(n924) );
    NAND2 U879 ( .O(n926), .I1(\mem<9><8> ), .I0(n322) );
    NAND2 U880 ( .O(n925), .I1(\mem<12><8> ), .I0(n325) );
    NAND2 U881 ( .O(n335), .I1(n925), .I0(n926) );
    NAND2 U882 ( .O(n928), .I1(\mem<10><8> ), .I0(n323) );
    NAND2 U883 ( .O(n927), .I1(\mem<13><8> ), .I0(n326) );
    NAND2 U884 ( .O(n334), .I1(n927), .I0(n928) );
    NAND2 U885 ( .O(n930), .I1(\mem<0><8> ), .I0(n314) );
    NAND2 U886 ( .O(n929), .I1(\mem<11><8> ), .I0(n324) );
    NAND2 U887 ( .O(n403), .I1(n929), .I0(n930) );
    NAND2 U888 ( .O(n932), .I1(\mem<1><8> ), .I0(n315) );
    NAND2 U889 ( .O(n931), .I1(n395), .I0(\mem<2><8> ) );
    NAND2 U890 ( .O(n402), .I1(n931), .I0(n932) );
    NAND2 U891 ( .O(n934), .I1(\mem<5><8> ), .I0(n317) );
    NAND2 U892 ( .O(n933), .I1(\mem<6><8> ), .I0(n318) );
    NAND2 U893 ( .O(n401), .I1(n933), .I0(n934) );
    NAND2 U894 ( .O(n936), .I1(\mem<4><8> ), .I0(n316) );
    NAND2 U895 ( .O(n935), .I1(n394), .I0(\mem<3><8> ) );
    NAND2 U896 ( .O(n400), .I1(n935), .I0(n936) );
    NAND2 U897 ( .O(n938), .I1(\mem<7><9> ), .I0(n319) );
    NAND2 U898 ( .O(n937), .I1(\mem<8><9> ), .I0(n321) );
    NAND2 U899 ( .O(n332), .I1(n937), .I0(n938) );
    NAND2 U900 ( .O(n940), .I1(\mem<9><9> ), .I0(n322) );
    NAND2 U901 ( .O(n939), .I1(\mem<12><9> ), .I0(n325) );
    NAND2 U902 ( .O(n331), .I1(n939), .I0(n940) );
    NAND2 U903 ( .O(n942), .I1(\mem<10><9> ), .I0(n323) );
    NAND2 U904 ( .O(n941), .I1(\mem<13><9> ), .I0(n326) );
    NAND2 U905 ( .O(n330), .I1(n941), .I0(n942) );
    NAND2 U906 ( .O(n944), .I1(\mem<0><9> ), .I0(n314) );
    NAND2 U907 ( .O(n943), .I1(\mem<11><9> ), .I0(n324) );
    NAND2 U908 ( .O(n399), .I1(n943), .I0(n944) );
    NAND2 U909 ( .O(n946), .I1(\mem<1><9> ), .I0(n315) );
    NAND2 U910 ( .O(n945), .I1(n395), .I0(\mem<2><9> ) );
    NAND2 U911 ( .O(n398), .I1(n945), .I0(n946) );
    NAND2 U912 ( .O(n948), .I1(\mem<5><9> ), .I0(n317) );
    NAND2 U913 ( .O(n947), .I1(\mem<6><9> ), .I0(n318) );
    NAND2 U914 ( .O(n397), .I1(n947), .I0(n948) );
    NAND2 U915 ( .O(n950), .I1(\mem<4><9> ), .I0(n316) );
    NAND2 U916 ( .O(n949), .I1(n394), .I0(\mem<3><9> ) );
    NAND2 U917 ( .O(n396), .I1(n949), .I0(n950) );
    INV U918 ( .O(n951), .I(n313) );
    INV U919 ( .O(n952), .I(n_14) );
    NOR4 U920 ( .O(n395), .I3(n_13), .I2(n_15), .I1(n951), .I0(n952) );
    INV U921 ( .O(n953), .I(n_13) );
    AND4 U922 ( .O(n394), .I3(n953), .I2(n313), .I1(n_14), .I0(n_15) );
    INV U923 ( .O(n955), .I(n954) );
    NAND2 U924 ( .O(n954), .I1(n147), .I0(n145) );
    OR2 U925 ( .O(\n68<0> ), .I1(\n55<9><9> ), .I0(n955) );
    INV U926 ( .O(n956), .I(n_12) );
    NOR3 U927 ( .O(n320), .I2(n_11), .I1(n_10), .I0(n956) );
    NOR3 U928 ( .O(n313), .I2(n_11), .I1(n_10), .I0(n_12) );
    INV U929 ( .O(n957), .I(n_14) );
    AND4 U930 ( .O(n326), .I3(n957), .I2(n320), .I1(n_15), .I0(n_13) );
    INV U931 ( .O(n958), .I(n320) );
    INV U932 ( .O(n959), .I(n_13) );
    NOR4 U933 ( .O(n325), .I3(n_15), .I2(n_14), .I1(n958), .I0(n959) );
    INV U934 ( .O(n960), .I(n_13) );
    AND4 U935 ( .O(n324), .I3(n960), .I2(n320), .I1(n_14), .I0(n_15) );
    INV U936 ( .O(n961), .I(n320) );
    INV U937 ( .O(n962), .I(n_14) );
    NOR4 U938 ( .O(n323), .I3(n_13), .I2(n_15), .I1(n961), .I0(n962) );
    INV U939 ( .O(n963), .I(n320) );
    INV U940 ( .O(n964), .I(n_15) );
    NOR4 U941 ( .O(n322), .I3(n_13), .I2(n_14), .I1(n963), .I0(n964) );
    INV U942 ( .O(n965), .I(n320) );
    NOR4 U943 ( .O(n321), .I3(n965), .I2(n_14), .I1(n_15), .I0(n_13) );
    AND4 U944 ( .O(n319), .I3(n313), .I2(n_14), .I1(n_15), .I0(n_13) );
    INV U945 ( .O(n966), .I(n_15) );
    AND4 U946 ( .O(n318), .I3(n966), .I2(n313), .I1(n_14), .I0(n_13) );
    INV U947 ( .O(n967), .I(n_14) );
    AND4 U948 ( .O(n317), .I3(n967), .I2(n313), .I1(n_15), .I0(n_13) );
    INV U949 ( .O(n968), .I(n313) );
    INV U950 ( .O(n969), .I(n_13) );
    NOR4 U951 ( .O(n316), .I3(n_15), .I2(n_14), .I1(n968), .I0(n969) );
    INV U952 ( .O(n970), .I(n313) );
    INV U953 ( .O(n971), .I(n_15) );
    NOR4 U954 ( .O(n315), .I3(n_13), .I2(n_14), .I1(n970), .I0(n971) );
    INV U955 ( .O(n972), .I(n313) );
    NOR4 U956 ( .O(n314), .I3(n972), .I2(n_14), .I1(n_15), .I0(n_13) );
    OR2 U957 ( .O(n974), .I1(n976), .I0(\n55<9><9> ) );
    NAND2 U958 ( .O(n973), .I1(\n55<9><9> ), .I0(n1068) );
    NAND2 U959 ( .O(n977), .I1(n973), .I0(n974) );
    NOR4 U960 ( .O(n976), .I3(n393), .I2(n392), .I1(n391), .I0(n390) );
    FDCE \data_bus_reg<0>  ( .Q(n1068), .D(n977), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U962 ( .O(n979), .I1(n981), .I0(\n55<9><9> ) );
    NAND2 U963 ( .O(n978), .I1(\n55<9><9> ), .I0(n1058) );
    NAND2 U964 ( .O(n982), .I1(n978), .I0(n979) );
    NOR4 U965 ( .O(n981), .I3(n389), .I2(n388), .I1(n387), .I0(n386) );
    FDCE \data_bus_reg<10>  ( .Q(n1058), .D(n982), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U967 ( .O(n984), .I1(n986), .I0(\n55<9><9> ) );
    NAND2 U968 ( .O(n983), .I1(\n55<9><9> ), .I0(n1057) );
    NAND2 U969 ( .O(n987), .I1(n983), .I0(n984) );
    NOR4 U970 ( .O(n986), .I3(n385), .I2(n384), .I1(n383), .I0(n382) );
    FDCE \data_bus_reg<11>  ( .Q(n1057), .D(n987), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U972 ( .O(n989), .I1(n991), .I0(\n55<9><9> ) );
    NAND2 U973 ( .O(n988), .I1(\n55<9><9> ), .I0(n1056) );
    NAND2 U974 ( .O(n992), .I1(n988), .I0(n989) );
    NOR4 U975 ( .O(n991), .I3(n381), .I2(n380), .I1(n379), .I0(n378) );
    FDCE \data_bus_reg<12>  ( .Q(n1056), .D(n992), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U977 ( .O(n994), .I1(n996), .I0(\n55<9><9> ) );
    NAND2 U978 ( .O(n993), .I1(\n55<9><9> ), .I0(n1055) );
    NAND2 U979 ( .O(n997), .I1(n993), .I0(n994) );
    NOR4 U980 ( .O(n996), .I3(n377), .I2(n376), .I1(n375), .I0(n374) );
    FDCE \data_bus_reg<13>  ( .Q(n1055), .D(n997), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U982 ( .O(n999), .I1(n1001), .I0(\n55<9><9> ) );
    NAND2 U983 ( .O(n998), .I1(\n55<9><9> ), .I0(n1054) );
    NAND2 U984 ( .O(n1002), .I1(n998), .I0(n999) );
    NOR4 U985 ( .O(n1001), .I3(n373), .I2(n372), .I1(n371), .I0(n370) );
    FDCE \data_bus_reg<14>  ( .Q(n1054), .D(n1002), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U987 ( .O(n1004), .I1(n1006), .I0(\n55<9><9> ) );
    NAND2 U988 ( .O(n1003), .I1(\n55<9><9> ), .I0(n1053) );
    NAND2 U989 ( .O(n1007), .I1(n1003), .I0(n1004) );
    NOR4 U990 ( .O(n1006), .I3(n369), .I2(n368), .I1(n367), .I0(n366) );
    FDCE \data_bus_reg<15>  ( .Q(n1053), .D(n1007), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U992 ( .O(n1009), .I1(n1011), .I0(\n55<9><9> ) );
    NAND2 U993 ( .O(n1008), .I1(\n55<9><9> ), .I0(n1067) );
    NAND2 U994 ( .O(n1012), .I1(n1008), .I0(n1009) );
    NOR4 U995 ( .O(n1011), .I3(n365), .I2(n364), .I1(n363), .I0(n362) );
    FDCE \data_bus_reg<1>  ( .Q(n1067), .D(n1012), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U997 ( .O(n1014), .I1(n1016), .I0(\n55<9><9> ) );
    NAND2 U998 ( .O(n1013), .I1(\n55<9><9> ), .I0(n1066) );
    NAND2 U999 ( .O(n1017), .I1(n1013), .I0(n1014) );
    NOR4 U1000 ( .O(n1016), .I3(n361), .I2(n360), .I1(n359), .I0(n358) );
    FDCE \data_bus_reg<2>  ( .Q(n1066), .D(n1017), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1002 ( .O(n1019), .I1(n1021), .I0(\n55<9><9> ) );
    NAND2 U1003 ( .O(n1018), .I1(\n55<9><9> ), .I0(n1065) );
    NAND2 U1004 ( .O(n1022), .I1(n1018), .I0(n1019) );
    NOR4 U1005 ( .O(n1021), .I3(n357), .I2(n356), .I1(n355), .I0(n354) );
    FDCE \data_bus_reg<3>  ( .Q(n1065), .D(n1022), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1007 ( .O(n1024), .I1(n1026), .I0(\n55<9><9> ) );
    NAND2 U1008 ( .O(n1023), .I1(\n55<9><9> ), .I0(n1064) );
    NAND2 U1009 ( .O(n1027), .I1(n1023), .I0(n1024) );
    NOR4 U1010 ( .O(n1026), .I3(n353), .I2(n352), .I1(n351), .I0(n350) );
    FDCE \data_bus_reg<4>  ( .Q(n1064), .D(n1027), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1012 ( .O(n1029), .I1(n1031), .I0(\n55<9><9> ) );
    NAND2 U1013 ( .O(n1028), .I1(\n55<9><9> ), .I0(n1063) );
    NAND2 U1014 ( .O(n1032), .I1(n1028), .I0(n1029) );
    NOR4 U1015 ( .O(n1031), .I3(n349), .I2(n348), .I1(n347), .I0(n346) );
    FDCE \data_bus_reg<5>  ( .Q(n1063), .D(n1032), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1017 ( .O(n1034), .I1(n1036), .I0(\n55<9><9> ) );
    NAND2 U1018 ( .O(n1033), .I1(\n55<9><9> ), .I0(n1062) );
    NAND2 U1019 ( .O(n1037), .I1(n1033), .I0(n1034) );
    NOR4 U1020 ( .O(n1036), .I3(n345), .I2(n344), .I1(n343), .I0(n342) );
    FDCE \data_bus_reg<6>  ( .Q(n1062), .D(n1037), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1022 ( .O(n1039), .I1(n1041), .I0(\n55<9><9> ) );
    NAND2 U1023 ( .O(n1038), .I1(\n55<9><9> ), .I0(n1061) );
    NAND2 U1024 ( .O(n1042), .I1(n1038), .I0(n1039) );
    NOR4 U1025 ( .O(n1041), .I3(n341), .I2(n340), .I1(n339), .I0(n338) );
    FDCE \data_bus_reg<7>  ( .Q(n1061), .D(n1042), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1027 ( .O(n1044), .I1(n1046), .I0(\n55<9><9> ) );
    NAND2 U1028 ( .O(n1043), .I1(\n55<9><9> ), .I0(n1060) );
    NAND2 U1029 ( .O(n1047), .I1(n1043), .I0(n1044) );
    NOR4 U1030 ( .O(n1046), .I3(n337), .I2(n336), .I1(n335), .I0(n334) );
    FDCE \data_bus_reg<8>  ( .Q(n1060), .D(n1047), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
    OR2 U1032 ( .O(n1049), .I1(n1051), .I0(\n55<9><9> ) );
    NAND2 U1033 ( .O(n1048), .I1(\n55<9><9> ), .I0(n1059) );
    NAND2 U1034 ( .O(n1052), .I1(n1048), .I0(n1049) );
    NOR4 U1035 ( .O(n1051), .I3(n333), .I2(n332), .I1(n331), .I0(n330) );
    FDCE \data_bus_reg<9>  ( .Q(n1059), .D(n1052), .C(n146), .CE(\n68<0> ), 
        .CLR(1'b0) );
endmodule

