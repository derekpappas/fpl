// Test type: Continuous assignment - pl1, st0 - list_of_net_assignments - 3 elements
// Vparser rule name:
// Author: andreib
module continuous393;
wire a,b,c;
assign (pull1, strong0) a=1'b1, b=1'b0, c=1'd2;
endmodule
