// Test type: loop statement - forever
// Vparser rule name:
// Author: andreib
module loop_statement1;
reg a;
initial forever a=1'b1;
endmodule
