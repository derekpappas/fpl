`include "defines.v"

module g0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 39
  input [1 - 1:0] ar_sa0_s10;
  f0 f0(.ar_sa0_s10(ar_sa0_s10));
  `include "g0.logic.vh"
endmodule

