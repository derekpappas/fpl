module Top_tb  ; 
 
  Top  
   DUT  ( ); 

endmodule

