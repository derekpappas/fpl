//test type : block_item_declaration ::= reg[signed][range] list_of_block_variable_identifiers;
//vparser rule name : 
//author : Codrin
module test_0480;
  (* sign = 1, regs *)
  reg signed [31:0] int1, int2, result;
endmodule
