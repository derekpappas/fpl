--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : b.vh
--FILE GENERATED ON : Sun Mar  7 15:39:23 2010

a.vhd
b.vhd
stim_expect_mem_template.vhd
tb.vhd
