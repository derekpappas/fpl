//test type : block_item_declaration ::= real list_of_block_variable_identifiers;
//vparser rule name : 
//author : Codrin
module test_0520;
  (* reset *)
  real value, result[1:10], exp;
endmodule
