`include "defines.v"

module u0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 143
  input [1 - 1:0] ar_sa0_s10;
  t0 t0(.ar_sa0_s10(ar_sa0_s10));
  `include "u0.logic.vh"
endmodule

