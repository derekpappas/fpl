// Test type: case_statement - case - 2 x expression:null
// Vparser rule name:
// Author: andreib
module case_statement11;
reg a;
initial case(a)
	4'b0000:;
	4'b0001:;
	endcase
endmodule
