//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : eth_mac.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module eth_mac(eb_emdummy4);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 26
  input eb_emdummy4;
  `include "eth_mac.logic.v"
endmodule

