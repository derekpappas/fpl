`include "defines.v"

module b_a1(x);
// Location of source csl unit: file name = gen_uniq_rtl1.csl line number = 15
  input x;
  `include "b_a1.logic.v"
endmodule

