localmem.vhd
localmem_register_file_memory.vhd
ctrlstore.vhd
execu.vhd
rf128.vhd
rf128_register_file_memory.vhd
crc.vhd
crcr.vhd
opmux.vhd
rfmux.vhd
msf.vhd
sramctrl.vhd
dramctrl.vhd
hash.vhd
pcictrl.vhd
cap.vhd
me.vhd
mecluster.vhd
xpi.vhd
dram.vhd
dram_register_file_memory.vhd
xscalecore.vhd
chip.vhd
