// Test type: Hex Numbers - 1 number
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=4'h3;
endmodule
