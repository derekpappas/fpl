-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./utop_cslc_generated/code/vhdl/u11.vhd
-- FILE GENERATED ON : Sat Mar 14 19:03:19 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u11\ is
  port(\ifcrc1_reset\ : in csl_bit;
       \ifcrc1_clock\ : in csl_bit;
       \ifc11_i0_pin\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \ifc11_i0_pout\ : out csl_bit_vector(10#8# - 10#1# downto 10#0#));
begin
end entity;

architecture \u11_logic\ of \u11\ is
begin
end architecture;

