`celldefine
module x;
endmodule

module y;
endmodule

module z;
endmodule
`endcelldefine


