//test type : port_declaration
//vparser rule name : 
//author : Codrin
module declaration_0130(x);
 (* a *) inout x;
endmodule
