// Test type: conditional_statement - if(expr) statement
// Vparser rule name:
// Author: andreib
module conditional_statement2;
reg a,b,c;
initial if(a==b) c=1;
endmodule
