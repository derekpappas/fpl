u1.vhd
u2.vhd
u3.vhd
u4.vhd
