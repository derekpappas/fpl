// Test type: Real numbers - exponent upper case sign
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=12.3E+12;
endmodule
