--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : top.vh
--FILE GENERATED ON : Thu Jun 10 02:45:25 2010

a.vhd
b.vhd
c.vhd
top.vhd
stim_expect_mem_template.vhd
tb.vhd
