// Test type: Real numbers - real number with underscore
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=27_4_.3_2_;
endmodule
