// Test type: Continuous assignment - sup1, st0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous271;
wire a;
assign (supply1, strong0) a=1'b1;
endmodule
