`include "defines.v"

module f1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 213
  output [1 - 1:0] ar_sa0_s10;
  e1 e10(.ar_sa0_s10(ar_sa0_s10));
  `include "f1.logic.vh"
endmodule

