// Test type: Real numbers - simple real exponential number
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1.3e9;
endmodule
