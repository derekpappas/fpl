`include "defines.v"

module e0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 25
  input [1 - 1:0] ar_sa0_s10;
  d0 d0(.ar_sa0_s10(ar_sa0_s10));
  `include "e0.logic.vh"
endmodule

