-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./ar15a_cslc_generated/code/vhdl/ud.vhd
-- FILE GENERATED ON : Sat Mar 14 17:54:45 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \ud\ is
  port(\pdin\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \pdout1\ : out csl_bit_vector(10#16# - 10#1# downto 10#0#);
       \pdout2\ : out csl_bit_vector(10#3# - 10#1# downto 10#0#);
       \ifcin_hw\ : in csl_bit_vector(10#16# - 10#1# downto 10#0#);
       \ifcin_w\ : in csl_bit_vector(10#8# - 10#1# downto 10#0#);
       \ifcrc_reset\ : in csl_bit;
       \ifcrc_clock\ : in csl_bit);
begin
end entity;

architecture \ud_logic\ of \ud\ is
begin
end architecture;

