-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./chip_cslc_generated/code/vhdl/u_rf.vhd
-- FILE GENERATED ON : Wed Nov 18 19:49:18 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_rf\ is
  port(\ifc_rf_p_clk\ : in csl_bit;
       \ifc_rf_p_rst\ : in csl_bit;
       \ifc_rf_p_stall\ : in csl_bit;
       \ifc_unit_rf_l_p_unitOut\ : out csl_bit_vector(10#32# - 10#1# downto 10#0#);
       \ifc_unit_rf_l_p_unitIn\ : in csl_bit_vector(10#32# - 10#1# downto 10#0#);
       \ifc_unit_rf_r_p_unitOut\ : out csl_bit_vector(10#32# - 10#1# downto 10#0#);
       \ifc_unit_rf_r_p_unitIn\ : in csl_bit_vector(10#32# - 10#1# downto 10#0#));
begin
end entity;

architecture \u_rf_logic\ of \u_rf\ is
begin
end architecture;

