// Test type: case_statement - case - expression:null
// Vparser rule name:
// Author: andreib
module case_statement1;
reg a;
initial case(a)
	4'b0000:;
	endcase
endmodule
