// Xilinx Verilog produced by program ngd2ver, Version M1.3.7
// Date: Wed Aug 13 17:58:11 1997
// Design file: /var/tmp/shifter_16.ngd
// Device: xc4000e
`timescale 1 ns/1 ps

  module shifter_16 (MS_IN, SYNC_CTRL, CLK_EN, CLOCK, Q_OUT);
    input MS_IN;
    input SYNC_CTRL;
    input CLK_EN;
    input CLOCK;
    output [15:0] Q_OUT;

    wire LB_GND, AND10_OUT, INV0_OUT, AND20_OUT, OR0_OUT, AND11_OUT, INV1_OUT, 
    AND21_OUT, OR1_OUT, AND12_OUT, INV2_OUT, AND22_OUT, OR2_OUT, AND13_OUT, 
    INV3_OUT, AND23_OUT, OR3_OUT, AND14_OUT, INV4_OUT, AND24_OUT, OR4_OUT, 
    AND15_OUT, INV5_OUT, AND25_OUT, OR5_OUT, AND16_OUT, INV6_OUT, AND26_OUT, 
    OR6_OUT, AND17_OUT, INV7_OUT, AND27_OUT, OR7_OUT, AND18_OUT, INV8_OUT, 
    AND28_OUT, OR8_OUT, AND19_OUT, INV9_OUT, AND29_OUT, OR9_OUT, AND110_OUT, 
    INV10_OUT, AND210_OUT, OR10_OUT, AND111_OUT, INV11_OUT, AND211_OUT, OR11_OUT
    , AND112_OUT, INV12_OUT, AND212_OUT, OR12_OUT, AND113_OUT, INV13_OUT, 
    AND213_OUT, OR13_OUT, AND114_OUT, INV14_OUT, AND214_OUT, OR14_OUT, 
    AND115_OUT, INV15_OUT, AND215_OUT, OR15_OUT, GND;
    `ifdef GSR_SIGNAL
      wire GSR = `GSR_SIGNAL ;
    `else
      wire GSR ;
    `endif

    X_ZERO LOGIC0 (.OUT (LB_GND));
    X_AND2 AND10 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND10_OUT));
    X_INV INV0 (.IN (SYNC_CTRL), .OUT (INV0_OUT));
    X_AND2 AND20 (.IN0 (Q_OUT[1]), .IN1 (INV0_OUT), .OUT (AND20_OUT));
    X_OR2 OR0 (.IN0 (AND10_OUT), .IN1 (AND20_OUT), .OUT (OR0_OUT));
    X_FF FF0 (.IN (OR0_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[0]));
    X_AND2 AND11 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND11_OUT));
    X_INV INV1 (.IN (SYNC_CTRL), .OUT (INV1_OUT));
    X_AND2 AND21 (.IN0 (Q_OUT[2]), .IN1 (INV1_OUT), .OUT (AND21_OUT));
    X_OR2 OR1 (.IN0 (AND11_OUT), .IN1 (AND21_OUT), .OUT (OR1_OUT));
    X_FF FF1 (.IN (OR1_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[1]));
    X_AND2 AND12 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND12_OUT));
    X_INV INV2 (.IN (SYNC_CTRL), .OUT (INV2_OUT));
    X_AND2 AND22 (.IN0 (Q_OUT[3]), .IN1 (INV2_OUT), .OUT (AND22_OUT));
    X_OR2 OR2 (.IN0 (AND12_OUT), .IN1 (AND22_OUT), .OUT (OR2_OUT));
    X_FF FF2 (.IN (OR2_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[2]));
    X_AND2 AND13 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND13_OUT));
    X_INV INV3 (.IN (SYNC_CTRL), .OUT (INV3_OUT));
    X_AND2 AND23 (.IN0 (Q_OUT[4]), .IN1 (INV3_OUT), .OUT (AND23_OUT));
    X_OR2 OR3 (.IN0 (AND13_OUT), .IN1 (AND23_OUT), .OUT (OR3_OUT));
    X_FF FF3 (.IN (OR3_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[3]));
    X_AND2 AND14 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND14_OUT));
    X_INV INV4 (.IN (SYNC_CTRL), .OUT (INV4_OUT));
    X_AND2 AND24 (.IN0 (Q_OUT[5]), .IN1 (INV4_OUT), .OUT (AND24_OUT));
    X_OR2 OR4 (.IN0 (AND14_OUT), .IN1 (AND24_OUT), .OUT (OR4_OUT));
    X_FF FF4 (.IN (OR4_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[4]));
    X_AND2 AND15 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND15_OUT));
    X_INV INV5 (.IN (SYNC_CTRL), .OUT (INV5_OUT));
    X_AND2 AND25 (.IN0 (Q_OUT[6]), .IN1 (INV5_OUT), .OUT (AND25_OUT));
    X_OR2 OR5 (.IN0 (AND15_OUT), .IN1 (AND25_OUT), .OUT (OR5_OUT));
    X_FF FF5 (.IN (OR5_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[5]));
    X_AND2 AND16 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND16_OUT));
    X_INV INV6 (.IN (SYNC_CTRL), .OUT (INV6_OUT));
    X_AND2 AND26 (.IN0 (Q_OUT[7]), .IN1 (INV6_OUT), .OUT (AND26_OUT));
    X_OR2 OR6 (.IN0 (AND16_OUT), .IN1 (AND26_OUT), .OUT (OR6_OUT));
    X_FF FF6 (.IN (OR6_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[6]));
    X_AND2 AND17 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND17_OUT));
    X_INV INV7 (.IN (SYNC_CTRL), .OUT (INV7_OUT));
    X_AND2 AND27 (.IN0 (Q_OUT[8]), .IN1 (INV7_OUT), .OUT (AND27_OUT));
    X_OR2 OR7 (.IN0 (AND17_OUT), .IN1 (AND27_OUT), .OUT (OR7_OUT));
    X_FF FF7 (.IN (OR7_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[7]));
    X_AND2 AND18 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND18_OUT));
    X_INV INV8 (.IN (SYNC_CTRL), .OUT (INV8_OUT));
    X_AND2 AND28 (.IN0 (Q_OUT[9]), .IN1 (INV8_OUT), .OUT (AND28_OUT));
    X_OR2 OR8 (.IN0 (AND18_OUT), .IN1 (AND28_OUT), .OUT (OR8_OUT));
    X_FF FF8 (.IN (OR8_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[8]));
    X_AND2 AND19 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND19_OUT));
    X_INV INV9 (.IN (SYNC_CTRL), .OUT (INV9_OUT));
    X_AND2 AND29 (.IN0 (Q_OUT[10]), .IN1 (INV9_OUT), .OUT (AND29_OUT));
    X_OR2 OR9 (.IN0 (AND19_OUT), .IN1 (AND29_OUT), .OUT (OR9_OUT));
    X_FF FF9 (.IN (OR9_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), .RST (GSR)
    , .OUT (Q_OUT[9]));
    X_AND2 AND110 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND110_OUT));
    X_INV INV10 (.IN (SYNC_CTRL), .OUT (INV10_OUT));
    X_AND2 AND210 (.IN0 (Q_OUT[11]), .IN1 (INV10_OUT), .OUT (AND210_OUT));
    X_OR2 OR10 (.IN0 (AND110_OUT), .IN1 (AND210_OUT), .OUT (OR10_OUT));
    X_FF FF10 (.IN (OR10_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), 
    .RST (GSR), .OUT (Q_OUT[10]));
    X_AND2 AND111 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND111_OUT));
    X_INV INV11 (.IN (SYNC_CTRL), .OUT (INV11_OUT));
    X_AND2 AND211 (.IN0 (Q_OUT[12]), .IN1 (INV11_OUT), .OUT (AND211_OUT));
    X_OR2 OR11 (.IN0 (AND111_OUT), .IN1 (AND211_OUT), .OUT (OR11_OUT));
    X_FF FF11 (.IN (OR11_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), 
    .RST (GSR), .OUT (Q_OUT[11]));
    X_AND2 AND112 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND112_OUT));
    X_INV INV12 (.IN (SYNC_CTRL), .OUT (INV12_OUT));
    X_AND2 AND212 (.IN0 (Q_OUT[13]), .IN1 (INV12_OUT), .OUT (AND212_OUT));
    X_OR2 OR12 (.IN0 (AND112_OUT), .IN1 (AND212_OUT), .OUT (OR12_OUT));
    X_FF FF12 (.IN (OR12_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), 
    .RST (GSR), .OUT (Q_OUT[12]));
    X_AND2 AND113 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND113_OUT));
    X_INV INV13 (.IN (SYNC_CTRL), .OUT (INV13_OUT));
    X_AND2 AND213 (.IN0 (Q_OUT[14]), .IN1 (INV13_OUT), .OUT (AND213_OUT));
    X_OR2 OR13 (.IN0 (AND113_OUT), .IN1 (AND213_OUT), .OUT (OR13_OUT));
    X_FF FF13 (.IN (OR13_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), 
    .RST (GSR), .OUT (Q_OUT[13]));
    X_AND2 AND114 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND114_OUT));
    X_INV INV14 (.IN (SYNC_CTRL), .OUT (INV14_OUT));
    X_AND2 AND214 (.IN0 (Q_OUT[15]), .IN1 (INV14_OUT), .OUT (AND214_OUT));
    X_OR2 OR14 (.IN0 (AND114_OUT), .IN1 (AND214_OUT), .OUT (OR14_OUT));
    X_FF FF14 (.IN (OR14_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), 
    .RST (GSR), .OUT (Q_OUT[14]));
    X_AND2 AND115 (.IN0 (LB_GND), .IN1 (SYNC_CTRL), .OUT (AND115_OUT));
    X_INV INV15 (.IN (SYNC_CTRL), .OUT (INV15_OUT));
    X_AND2 AND215 (.IN0 (MS_IN), .IN1 (INV15_OUT), .OUT (AND215_OUT));
    X_OR2 OR15 (.IN0 (AND115_OUT), .IN1 (AND215_OUT), .OUT (OR15_OUT));
    X_FF FF15 (.IN (OR15_OUT), .CLK (CLOCK), .CE (CLK_EN), .SET (GND), 
    .RST (GSR), .OUT (Q_OUT[15]));
    X_ZERO GND_82 (.OUT (GND));
    X_PD NGD2VER_PD_85 (.OUT (GSR) );
  endmodule

