// Test type: Decimal Numbers - 0 preceded decimal number
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=023;
endmodule
