-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./b_cslc_generated/code/vhdl/a.vhd
-- FILE GENERATED ON : Mon Nov 16 08:40:43 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \a\ is
  port(\in_a\ : in csl_bit;
       \out_a\ : out csl_bit;
       \clk\ : in csl_bit);
begin
end entity;

architecture \a_logic\ of \a\ is
begin
end architecture;

