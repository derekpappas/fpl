//test type : task_item_declaration ::= output_declaration
//vparser rule name : 
//author : Codrin
//fixed by: Gabrield
module test_0460;
 task add(
  (* cout, cin *)
  output sum);
  ;
 endtask
endmodule
