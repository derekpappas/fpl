// Test type: initial statement - procedural_continuous_assign - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon25;
reg [7:0]a;
initial 
assign a=2;
endmodule
