// Test type: Decimal Numbers - lower case signed upper case decimal base
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'sD2___9;
endmodule
