//test type : operator_~^ system_funtion_call
//vparser rule name : 
//author : Bogdan Mereghea
module unary_operator65;
    wire a;
    assign a = ~^$random;
endmodule
