//test type : module_or_generate_item ::= module_or_generate_item_declaration (realtime_declaration)
//vparser rule name : 
//author : Codrin
module test_0210;
 (* realtimed = 1, treal =0, rtime = 0 *) realtime rtime[1:6];
endmodule
