module testbench_reg_declaration;
    reg_declaration0 reg_declaration_instance0();
    reg_declaration1 reg_declaration_instance1();
    reg_declaration2 reg_declaration_instance2();
    reg_declaration3 reg_declaration_instance3();
    reg_declaration4 reg_declaration_instance4();
    reg_declaration5 reg_declaration_instance5();
    reg_declaration6 reg_declaration_instance6();
    reg_declaration7 reg_declaration_instance7();
    reg_declaration8 reg_declaration_instance8();
    reg_declaration9 reg_declaration_instance9();
    reg_declaration10 reg_declaration_instance10();
    reg_declaration11 reg_declaration_instance11();
    reg_declaration12 reg_declaration_instance12();
    reg_declaration13 reg_declaration_instance13();
    reg_declaration14 reg_declaration_instance14();
    reg_declaration15 reg_declaration_instance15();
    reg_declaration16 reg_declaration_instance16();
    reg_declaration17 reg_declaration_instance17();
    reg_declaration18 reg_declaration_instance18();
    reg_declaration19 reg_declaration_instance19();
    reg_declaration20 reg_declaration_instance20();
    reg_declaration21 reg_declaration_instance21();
    reg_declaration22 reg_declaration_instance22();
    reg_declaration23 reg_declaration_instance23();
    reg_declaration24 reg_declaration_instance24();
    reg_declaration25 reg_declaration_instance25();
    reg_declaration26 reg_declaration_instance26();
    reg_declaration27 reg_declaration_instance27();
    reg_declaration28 reg_declaration_instance28();
    reg_declaration29 reg_declaration_instance29();
    reg_declaration30 reg_declaration_instance30();
    reg_declaration31 reg_declaration_instance31();
    reg_declaration32 reg_declaration_instance32();
    reg_declaration33 reg_declaration_instance33();
    reg_declaration34 reg_declaration_instance34();
    reg_declaration35 reg_declaration_instance35();
    reg_declaration36 reg_declaration_instance36();
    reg_declaration37 reg_declaration_instance37();
    reg_declaration38 reg_declaration_instance38();
    reg_declaration39 reg_declaration_instance39();
    reg_declaration40 reg_declaration_instance40();
    reg_declaration41 reg_declaration_instance41();
    reg_declaration42 reg_declaration_instance42();
    reg_declaration43 reg_declaration_instance43();
    reg_declaration44 reg_declaration_instance44();
    reg_declaration45 reg_declaration_instance45();
    reg_declaration46 reg_declaration_instance46();
    reg_declaration47 reg_declaration_instance47();
    reg_declaration48 reg_declaration_instance48();
    reg_declaration49 reg_declaration_instance49();
    reg_declaration50 reg_declaration_instance50();
    reg_declaration51 reg_declaration_instance51();
    reg_declaration52 reg_declaration_instance52();
    reg_declaration53 reg_declaration_instance53();
    reg_declaration54 reg_declaration_instance54();
    reg_declaration55 reg_declaration_instance55();
    reg_declaration56 reg_declaration_instance56();
    reg_declaration57 reg_declaration_instance57();
    reg_declaration58 reg_declaration_instance58();
    reg_declaration59 reg_declaration_instance59();
    reg_declaration60 reg_declaration_instance60();
    reg_declaration61 reg_declaration_instance61();
    reg_declaration62 reg_declaration_instance62();
    reg_declaration63 reg_declaration_instance63();
    reg_declaration64 reg_declaration_instance64();
    reg_declaration65 reg_declaration_instance65();
    reg_declaration66 reg_declaration_instance66();
    reg_declaration67 reg_declaration_instance67();
    reg_declaration68 reg_declaration_instance68();
    reg_declaration69 reg_declaration_instance69();
    reg_declaration70 reg_declaration_instance70();
    reg_declaration71 reg_declaration_instance71();
    reg_declaration72 reg_declaration_instance72();
    reg_declaration73 reg_declaration_instance73();
    reg_declaration74 reg_declaration_instance74();
    reg_declaration75 reg_declaration_instance75();
    reg_declaration76 reg_declaration_instance76();
    reg_declaration77 reg_declaration_instance77();
    reg_declaration78 reg_declaration_instance78();
    reg_declaration79 reg_declaration_instance79();
    reg_declaration80 reg_declaration_instance80();
    reg_declaration81 reg_declaration_instance81();
    reg_declaration82 reg_declaration_instance82();
    reg_declaration83 reg_declaration_instance83();
    reg_declaration84 reg_declaration_instance84();
    reg_declaration85 reg_declaration_instance85();
    reg_declaration86 reg_declaration_instance86();
    reg_declaration87 reg_declaration_instance87();
    reg_declaration88 reg_declaration_instance88();
    reg_declaration89 reg_declaration_instance89();
    reg_declaration90 reg_declaration_instance90();
    reg_declaration91 reg_declaration_instance91();
    reg_declaration92 reg_declaration_instance92();
    reg_declaration93 reg_declaration_instance93();
    reg_declaration94 reg_declaration_instance94();
    reg_declaration95 reg_declaration_instance95();
    reg_declaration96 reg_declaration_instance96();
    reg_declaration97 reg_declaration_instance97();
    reg_declaration98 reg_declaration_instance98();
    reg_declaration99 reg_declaration_instance99();
    reg_declaration100 reg_declaration_instance100();
    reg_declaration101 reg_declaration_instance101();
    reg_declaration102 reg_declaration_instance102();
    reg_declaration103 reg_declaration_instance103();
    reg_declaration104 reg_declaration_instance104();
    reg_declaration105 reg_declaration_instance105();
    reg_declaration106 reg_declaration_instance106();
    reg_declaration107 reg_declaration_instance107();
    reg_declaration108 reg_declaration_instance108();
    reg_declaration109 reg_declaration_instance109();
    reg_declaration110 reg_declaration_instance110();
    reg_declaration111 reg_declaration_instance111();
    reg_declaration112 reg_declaration_instance112();
    reg_declaration113 reg_declaration_instance113();
    reg_declaration114 reg_declaration_instance114();
    reg_declaration115 reg_declaration_instance115();
    reg_declaration116 reg_declaration_instance116();
    reg_declaration117 reg_declaration_instance117();
    reg_declaration118 reg_declaration_instance118();
    reg_declaration119 reg_declaration_instance119();
    reg_declaration120 reg_declaration_instance120();
    reg_declaration121 reg_declaration_instance121();
    reg_declaration122 reg_declaration_instance122();
    reg_declaration123 reg_declaration_instance123();
    reg_declaration124 reg_declaration_instance124();
    reg_declaration125 reg_declaration_instance125();
    reg_declaration126 reg_declaration_instance126();
    reg_declaration127 reg_declaration_instance127();
    reg_declaration128 reg_declaration_instance128();
    reg_declaration129 reg_declaration_instance129();
    reg_declaration130 reg_declaration_instance130();
    reg_declaration131 reg_declaration_instance131();
    reg_declaration132 reg_declaration_instance132();
    reg_declaration133 reg_declaration_instance133();
    reg_declaration134 reg_declaration_instance134();
    reg_declaration135 reg_declaration_instance135();
    reg_declaration136 reg_declaration_instance136();
    reg_declaration137 reg_declaration_instance137();
    reg_declaration138 reg_declaration_instance138();
    reg_declaration139 reg_declaration_instance139();
    reg_declaration140 reg_declaration_instance140();
    reg_declaration141 reg_declaration_instance141();
    reg_declaration142 reg_declaration_instance142();
    reg_declaration143 reg_declaration_instance143();
    reg_declaration144 reg_declaration_instance144();
    reg_declaration145 reg_declaration_instance145();
    reg_declaration146 reg_declaration_instance146();
    reg_declaration147 reg_declaration_instance147();
    reg_declaration148 reg_declaration_instance148();
    reg_declaration149 reg_declaration_instance149();
    reg_declaration150 reg_declaration_instance150();
    reg_declaration151 reg_declaration_instance151();
    reg_declaration152 reg_declaration_instance152();
    reg_declaration153 reg_declaration_instance153();
    reg_declaration154 reg_declaration_instance154();
    reg_declaration155 reg_declaration_instance155();
    reg_declaration156 reg_declaration_instance156();
    reg_declaration157 reg_declaration_instance157();
    reg_declaration158 reg_declaration_instance158();
    reg_declaration159 reg_declaration_instance159();
    reg_declaration160 reg_declaration_instance160();
    reg_declaration161 reg_declaration_instance161();
    reg_declaration162 reg_declaration_instance162();
    reg_declaration163 reg_declaration_instance163();
    reg_declaration164 reg_declaration_instance164();
    reg_declaration165 reg_declaration_instance165();
    reg_declaration166 reg_declaration_instance166();
    reg_declaration167 reg_declaration_instance167();
    reg_declaration168 reg_declaration_instance168();
    reg_declaration169 reg_declaration_instance169();
    reg_declaration170 reg_declaration_instance170();
    reg_declaration171 reg_declaration_instance171();
    reg_declaration172 reg_declaration_instance172();
    reg_declaration173 reg_declaration_instance173();
    reg_declaration174 reg_declaration_instance174();
    reg_declaration175 reg_declaration_instance175();
    reg_declaration176 reg_declaration_instance176();
    reg_declaration177 reg_declaration_instance177();
    reg_declaration178 reg_declaration_instance178();
    reg_declaration179 reg_declaration_instance179();
    reg_declaration180 reg_declaration_instance180();
    reg_declaration181 reg_declaration_instance181();
    reg_declaration182 reg_declaration_instance182();
    reg_declaration183 reg_declaration_instance183();
    reg_declaration184 reg_declaration_instance184();
    reg_declaration185 reg_declaration_instance185();
    reg_declaration186 reg_declaration_instance186();
    reg_declaration187 reg_declaration_instance187();
    reg_declaration188 reg_declaration_instance188();
    reg_declaration189 reg_declaration_instance189();
    reg_declaration190 reg_declaration_instance190();
    reg_declaration191 reg_declaration_instance191();
    reg_declaration192 reg_declaration_instance192();
    reg_declaration193 reg_declaration_instance193();
    reg_declaration194 reg_declaration_instance194();
    reg_declaration195 reg_declaration_instance195();
    reg_declaration196 reg_declaration_instance196();
    reg_declaration197 reg_declaration_instance197();
    reg_declaration198 reg_declaration_instance198();
    reg_declaration199 reg_declaration_instance199();
    reg_declaration200 reg_declaration_instance200();
    reg_declaration201 reg_declaration_instance201();
    reg_declaration202 reg_declaration_instance202();
    reg_declaration203 reg_declaration_instance203();
    reg_declaration204 reg_declaration_instance204();
    reg_declaration205 reg_declaration_instance205();
    reg_declaration206 reg_declaration_instance206();
    reg_declaration207 reg_declaration_instance207();
    reg_declaration208 reg_declaration_instance208();
    reg_declaration209 reg_declaration_instance209();
    reg_declaration210 reg_declaration_instance210();
    reg_declaration211 reg_declaration_instance211();
    reg_declaration212 reg_declaration_instance212();
    reg_declaration213 reg_declaration_instance213();
    reg_declaration214 reg_declaration_instance214();
    reg_declaration215 reg_declaration_instance215();
    reg_declaration216 reg_declaration_instance216();
    reg_declaration217 reg_declaration_instance217();
    reg_declaration218 reg_declaration_instance218();
    reg_declaration219 reg_declaration_instance219();
    reg_declaration220 reg_declaration_instance220();
    reg_declaration221 reg_declaration_instance221();
    reg_declaration222 reg_declaration_instance222();
    reg_declaration223 reg_declaration_instance223();
    reg_declaration224 reg_declaration_instance224();
    reg_declaration225 reg_declaration_instance225();
    reg_declaration226 reg_declaration_instance226();
    reg_declaration227 reg_declaration_instance227();
    reg_declaration228 reg_declaration_instance228();
    reg_declaration229 reg_declaration_instance229();
    reg_declaration230 reg_declaration_instance230();
    reg_declaration231 reg_declaration_instance231();
    reg_declaration232 reg_declaration_instance232();
    reg_declaration233 reg_declaration_instance233();
    reg_declaration234 reg_declaration_instance234();
    reg_declaration235 reg_declaration_instance235();
    reg_declaration236 reg_declaration_instance236();
    reg_declaration237 reg_declaration_instance237();
    reg_declaration238 reg_declaration_instance238();
    reg_declaration239 reg_declaration_instance239();
    reg_declaration240 reg_declaration_instance240();
    reg_declaration241 reg_declaration_instance241();
    reg_declaration242 reg_declaration_instance242();
    reg_declaration243 reg_declaration_instance243();
    reg_declaration244 reg_declaration_instance244();
    reg_declaration245 reg_declaration_instance245();
    reg_declaration246 reg_declaration_instance246();
    reg_declaration247 reg_declaration_instance247();
    reg_declaration248 reg_declaration_instance248();
    reg_declaration249 reg_declaration_instance249();
    reg_declaration250 reg_declaration_instance250();
    reg_declaration251 reg_declaration_instance251();
    reg_declaration252 reg_declaration_instance252();
    reg_declaration253 reg_declaration_instance253();
    reg_declaration254 reg_declaration_instance254();
    reg_declaration255 reg_declaration_instance255();
    reg_declaration256 reg_declaration_instance256();
    reg_declaration257 reg_declaration_instance257();
    reg_declaration258 reg_declaration_instance258();
    reg_declaration259 reg_declaration_instance259();
    reg_declaration260 reg_declaration_instance260();
    reg_declaration261 reg_declaration_instance261();
    reg_declaration262 reg_declaration_instance262();
    reg_declaration263 reg_declaration_instance263();
    reg_declaration264 reg_declaration_instance264();
    reg_declaration265 reg_declaration_instance265();
    reg_declaration266 reg_declaration_instance266();
    reg_declaration267 reg_declaration_instance267();
    reg_declaration268 reg_declaration_instance268();
    reg_declaration269 reg_declaration_instance269();
    reg_declaration270 reg_declaration_instance270();
    reg_declaration271 reg_declaration_instance271();
    reg_declaration272 reg_declaration_instance272();
    reg_declaration273 reg_declaration_instance273();
    reg_declaration274 reg_declaration_instance274();
    reg_declaration275 reg_declaration_instance275();
    reg_declaration276 reg_declaration_instance276();
    reg_declaration277 reg_declaration_instance277();
    reg_declaration278 reg_declaration_instance278();
    reg_declaration279 reg_declaration_instance279();
    reg_declaration280 reg_declaration_instance280();
    reg_declaration281 reg_declaration_instance281();
    reg_declaration282 reg_declaration_instance282();
    reg_declaration283 reg_declaration_instance283();
    reg_declaration284 reg_declaration_instance284();
    reg_declaration285 reg_declaration_instance285();
    reg_declaration286 reg_declaration_instance286();
    reg_declaration287 reg_declaration_instance287();
    reg_declaration288 reg_declaration_instance288();
    reg_declaration289 reg_declaration_instance289();
    reg_declaration290 reg_declaration_instance290();
    reg_declaration291 reg_declaration_instance291();
    reg_declaration292 reg_declaration_instance292();
    reg_declaration293 reg_declaration_instance293();
    reg_declaration294 reg_declaration_instance294();
    reg_declaration295 reg_declaration_instance295();
    reg_declaration296 reg_declaration_instance296();
    reg_declaration297 reg_declaration_instance297();
    reg_declaration298 reg_declaration_instance298();
    reg_declaration299 reg_declaration_instance299();
    reg_declaration300 reg_declaration_instance300();
    reg_declaration301 reg_declaration_instance301();
    reg_declaration302 reg_declaration_instance302();
    reg_declaration303 reg_declaration_instance303();
    reg_declaration304 reg_declaration_instance304();
    reg_declaration305 reg_declaration_instance305();
    reg_declaration306 reg_declaration_instance306();
    reg_declaration307 reg_declaration_instance307();
    reg_declaration308 reg_declaration_instance308();
    reg_declaration309 reg_declaration_instance309();
    reg_declaration310 reg_declaration_instance310();
    reg_declaration311 reg_declaration_instance311();
    reg_declaration312 reg_declaration_instance312();
    reg_declaration313 reg_declaration_instance313();
    reg_declaration314 reg_declaration_instance314();
    reg_declaration315 reg_declaration_instance315();
    reg_declaration316 reg_declaration_instance316();
    reg_declaration317 reg_declaration_instance317();
    reg_declaration318 reg_declaration_instance318();
    reg_declaration319 reg_declaration_instance319();
    reg_declaration320 reg_declaration_instance320();
    reg_declaration321 reg_declaration_instance321();
    reg_declaration322 reg_declaration_instance322();
    reg_declaration323 reg_declaration_instance323();
    reg_declaration324 reg_declaration_instance324();
    reg_declaration325 reg_declaration_instance325();
    reg_declaration326 reg_declaration_instance326();
    reg_declaration327 reg_declaration_instance327();
    reg_declaration328 reg_declaration_instance328();
    reg_declaration329 reg_declaration_instance329();
    reg_declaration330 reg_declaration_instance330();
    reg_declaration331 reg_declaration_instance331();
    reg_declaration332 reg_declaration_instance332();
    reg_declaration333 reg_declaration_instance333();
    reg_declaration334 reg_declaration_instance334();
    reg_declaration335 reg_declaration_instance335();
    reg_declaration336 reg_declaration_instance336();
    reg_declaration337 reg_declaration_instance337();
    reg_declaration338 reg_declaration_instance338();
    reg_declaration339 reg_declaration_instance339();
    reg_declaration340 reg_declaration_instance340();
    reg_declaration341 reg_declaration_instance341();
    reg_declaration342 reg_declaration_instance342();
    reg_declaration343 reg_declaration_instance343();
    reg_declaration344 reg_declaration_instance344();
    reg_declaration345 reg_declaration_instance345();
    reg_declaration346 reg_declaration_instance346();
    reg_declaration347 reg_declaration_instance347();
    reg_declaration348 reg_declaration_instance348();
    reg_declaration349 reg_declaration_instance349();
    reg_declaration350 reg_declaration_instance350();
    reg_declaration351 reg_declaration_instance351();
    reg_declaration352 reg_declaration_instance352();
    reg_declaration353 reg_declaration_instance353();
    reg_declaration354 reg_declaration_instance354();
    reg_declaration355 reg_declaration_instance355();
    reg_declaration356 reg_declaration_instance356();
    reg_declaration357 reg_declaration_instance357();
    reg_declaration358 reg_declaration_instance358();
    reg_declaration359 reg_declaration_instance359();
    reg_declaration360 reg_declaration_instance360();
    reg_declaration361 reg_declaration_instance361();
    reg_declaration362 reg_declaration_instance362();
    reg_declaration363 reg_declaration_instance363();
    reg_declaration364 reg_declaration_instance364();
    reg_declaration365 reg_declaration_instance365();
    reg_declaration366 reg_declaration_instance366();
    reg_declaration367 reg_declaration_instance367();
    reg_declaration368 reg_declaration_instance368();
    reg_declaration369 reg_declaration_instance369();
    reg_declaration370 reg_declaration_instance370();
    reg_declaration371 reg_declaration_instance371();
    reg_declaration372 reg_declaration_instance372();
    reg_declaration373 reg_declaration_instance373();
    reg_declaration374 reg_declaration_instance374();
    reg_declaration375 reg_declaration_instance375();
    reg_declaration376 reg_declaration_instance376();
    reg_declaration377 reg_declaration_instance377();
    reg_declaration378 reg_declaration_instance378();
    reg_declaration379 reg_declaration_instance379();
    reg_declaration380 reg_declaration_instance380();
    reg_declaration381 reg_declaration_instance381();
    reg_declaration382 reg_declaration_instance382();
    reg_declaration383 reg_declaration_instance383();
    reg_declaration384 reg_declaration_instance384();
    reg_declaration385 reg_declaration_instance385();
    reg_declaration386 reg_declaration_instance386();
    reg_declaration387 reg_declaration_instance387();
    reg_declaration388 reg_declaration_instance388();
    reg_declaration389 reg_declaration_instance389();
    reg_declaration390 reg_declaration_instance390();
    reg_declaration391 reg_declaration_instance391();
    reg_declaration392 reg_declaration_instance392();
    reg_declaration393 reg_declaration_instance393();
    reg_declaration394 reg_declaration_instance394();
    reg_declaration395 reg_declaration_instance395();
    reg_declaration396 reg_declaration_instance396();
    reg_declaration397 reg_declaration_instance397();
    reg_declaration398 reg_declaration_instance398();
    reg_declaration399 reg_declaration_instance399();
    reg_declaration400 reg_declaration_instance400();
    reg_declaration401 reg_declaration_instance401();
    reg_declaration402 reg_declaration_instance402();
    reg_declaration403 reg_declaration_instance403();
    reg_declaration404 reg_declaration_instance404();
    reg_declaration405 reg_declaration_instance405();
    reg_declaration406 reg_declaration_instance406();
    reg_declaration407 reg_declaration_instance407();
    reg_declaration408 reg_declaration_instance408();
    reg_declaration409 reg_declaration_instance409();
    reg_declaration410 reg_declaration_instance410();
    reg_declaration411 reg_declaration_instance411();
    reg_declaration412 reg_declaration_instance412();
    reg_declaration413 reg_declaration_instance413();
    reg_declaration414 reg_declaration_instance414();
    reg_declaration415 reg_declaration_instance415();
    reg_declaration416 reg_declaration_instance416();
    reg_declaration417 reg_declaration_instance417();
    reg_declaration418 reg_declaration_instance418();
    reg_declaration419 reg_declaration_instance419();
    reg_declaration420 reg_declaration_instance420();
    reg_declaration421 reg_declaration_instance421();
    reg_declaration422 reg_declaration_instance422();
    reg_declaration423 reg_declaration_instance423();
    reg_declaration424 reg_declaration_instance424();
    reg_declaration425 reg_declaration_instance425();
    reg_declaration426 reg_declaration_instance426();
    reg_declaration427 reg_declaration_instance427();
    reg_declaration428 reg_declaration_instance428();
    reg_declaration429 reg_declaration_instance429();
    reg_declaration430 reg_declaration_instance430();
    reg_declaration431 reg_declaration_instance431();
    reg_declaration432 reg_declaration_instance432();
    reg_declaration433 reg_declaration_instance433();
    reg_declaration434 reg_declaration_instance434();
    reg_declaration435 reg_declaration_instance435();
    reg_declaration436 reg_declaration_instance436();
    reg_declaration437 reg_declaration_instance437();
    reg_declaration438 reg_declaration_instance438();
    reg_declaration439 reg_declaration_instance439();
    reg_declaration440 reg_declaration_instance440();
    reg_declaration441 reg_declaration_instance441();
    reg_declaration442 reg_declaration_instance442();
    reg_declaration443 reg_declaration_instance443();
    reg_declaration444 reg_declaration_instance444();
    reg_declaration445 reg_declaration_instance445();
    reg_declaration446 reg_declaration_instance446();
    reg_declaration447 reg_declaration_instance447();
    reg_declaration448 reg_declaration_instance448();
    reg_declaration449 reg_declaration_instance449();
    reg_declaration450 reg_declaration_instance450();
    reg_declaration451 reg_declaration_instance451();
    reg_declaration452 reg_declaration_instance452();
    reg_declaration453 reg_declaration_instance453();
    reg_declaration454 reg_declaration_instance454();
    reg_declaration455 reg_declaration_instance455();
    reg_declaration456 reg_declaration_instance456();
    reg_declaration457 reg_declaration_instance457();
    reg_declaration458 reg_declaration_instance458();
    reg_declaration459 reg_declaration_instance459();
    reg_declaration460 reg_declaration_instance460();
    reg_declaration461 reg_declaration_instance461();
    reg_declaration462 reg_declaration_instance462();
    reg_declaration463 reg_declaration_instance463();
    reg_declaration464 reg_declaration_instance464();
    reg_declaration465 reg_declaration_instance465();
    reg_declaration466 reg_declaration_instance466();
    reg_declaration467 reg_declaration_instance467();
    reg_declaration468 reg_declaration_instance468();
    reg_declaration469 reg_declaration_instance469();
    reg_declaration470 reg_declaration_instance470();
    reg_declaration471 reg_declaration_instance471();
    reg_declaration472 reg_declaration_instance472();
    reg_declaration473 reg_declaration_instance473();
    reg_declaration474 reg_declaration_instance474();
    reg_declaration475 reg_declaration_instance475();
    reg_declaration476 reg_declaration_instance476();
    reg_declaration477 reg_declaration_instance477();
    reg_declaration478 reg_declaration_instance478();
    reg_declaration479 reg_declaration_instance479();
    reg_declaration480 reg_declaration_instance480();
    reg_declaration481 reg_declaration_instance481();
    reg_declaration482 reg_declaration_instance482();
    reg_declaration483 reg_declaration_instance483();
    reg_declaration484 reg_declaration_instance484();
    reg_declaration485 reg_declaration_instance485();
    reg_declaration486 reg_declaration_instance486();
    reg_declaration487 reg_declaration_instance487();
    reg_declaration488 reg_declaration_instance488();
    reg_declaration489 reg_declaration_instance489();
    reg_declaration490 reg_declaration_instance490();
    reg_declaration491 reg_declaration_instance491();
    reg_declaration492 reg_declaration_instance492();
    reg_declaration493 reg_declaration_instance493();
    reg_declaration494 reg_declaration_instance494();
    reg_declaration495 reg_declaration_instance495();
    reg_declaration496 reg_declaration_instance496();
    reg_declaration497 reg_declaration_instance497();
    reg_declaration498 reg_declaration_instance498();
    reg_declaration499 reg_declaration_instance499();
    reg_declaration500 reg_declaration_instance500();
    reg_declaration501 reg_declaration_instance501();
    reg_declaration502 reg_declaration_instance502();
    reg_declaration503 reg_declaration_instance503();
    reg_declaration504 reg_declaration_instance504();
    reg_declaration505 reg_declaration_instance505();
    reg_declaration506 reg_declaration_instance506();
    reg_declaration507 reg_declaration_instance507();
    reg_declaration508 reg_declaration_instance508();
    reg_declaration509 reg_declaration_instance509();
    reg_declaration510 reg_declaration_instance510();
    reg_declaration511 reg_declaration_instance511();
    reg_declaration512 reg_declaration_instance512();
    reg_declaration513 reg_declaration_instance513();
    reg_declaration514 reg_declaration_instance514();
    reg_declaration515 reg_declaration_instance515();
    reg_declaration516 reg_declaration_instance516();
    reg_declaration517 reg_declaration_instance517();
    reg_declaration518 reg_declaration_instance518();
    reg_declaration519 reg_declaration_instance519();
    reg_declaration520 reg_declaration_instance520();
    reg_declaration521 reg_declaration_instance521();
    reg_declaration522 reg_declaration_instance522();
    reg_declaration523 reg_declaration_instance523();
    reg_declaration524 reg_declaration_instance524();
    reg_declaration525 reg_declaration_instance525();
    reg_declaration526 reg_declaration_instance526();
    reg_declaration527 reg_declaration_instance527();
    reg_declaration528 reg_declaration_instance528();
    reg_declaration529 reg_declaration_instance529();
    reg_declaration530 reg_declaration_instance530();
    reg_declaration531 reg_declaration_instance531();
    reg_declaration532 reg_declaration_instance532();
    reg_declaration533 reg_declaration_instance533();
    reg_declaration534 reg_declaration_instance534();
    reg_declaration535 reg_declaration_instance535();
    reg_declaration536 reg_declaration_instance536();
    reg_declaration537 reg_declaration_instance537();
    reg_declaration538 reg_declaration_instance538();
    reg_declaration539 reg_declaration_instance539();
    reg_declaration540 reg_declaration_instance540();
    reg_declaration541 reg_declaration_instance541();
    reg_declaration542 reg_declaration_instance542();
    reg_declaration543 reg_declaration_instance543();
    reg_declaration544 reg_declaration_instance544();
    reg_declaration545 reg_declaration_instance545();
    reg_declaration546 reg_declaration_instance546();
    reg_declaration547 reg_declaration_instance547();
    reg_declaration548 reg_declaration_instance548();
    reg_declaration549 reg_declaration_instance549();
    reg_declaration550 reg_declaration_instance550();
    reg_declaration551 reg_declaration_instance551();
    reg_declaration552 reg_declaration_instance552();
    reg_declaration553 reg_declaration_instance553();
    reg_declaration554 reg_declaration_instance554();
    reg_declaration555 reg_declaration_instance555();
    reg_declaration556 reg_declaration_instance556();
    reg_declaration557 reg_declaration_instance557();
    reg_declaration558 reg_declaration_instance558();
    reg_declaration559 reg_declaration_instance559();
    reg_declaration560 reg_declaration_instance560();
    reg_declaration561 reg_declaration_instance561();
    reg_declaration562 reg_declaration_instance562();
    reg_declaration563 reg_declaration_instance563();
    reg_declaration564 reg_declaration_instance564();
    reg_declaration565 reg_declaration_instance565();
    reg_declaration566 reg_declaration_instance566();
    reg_declaration567 reg_declaration_instance567();
    reg_declaration568 reg_declaration_instance568();
    reg_declaration569 reg_declaration_instance569();
    reg_declaration570 reg_declaration_instance570();
    reg_declaration571 reg_declaration_instance571();
    reg_declaration572 reg_declaration_instance572();
    reg_declaration573 reg_declaration_instance573();
    reg_declaration574 reg_declaration_instance574();
    reg_declaration575 reg_declaration_instance575();
    reg_declaration576 reg_declaration_instance576();
    reg_declaration577 reg_declaration_instance577();
    reg_declaration578 reg_declaration_instance578();
    reg_declaration579 reg_declaration_instance579();
    reg_declaration580 reg_declaration_instance580();
    reg_declaration581 reg_declaration_instance581();
    reg_declaration582 reg_declaration_instance582();
    reg_declaration583 reg_declaration_instance583();
    reg_declaration584 reg_declaration_instance584();
    reg_declaration585 reg_declaration_instance585();
    reg_declaration586 reg_declaration_instance586();
    reg_declaration587 reg_declaration_instance587();
    reg_declaration588 reg_declaration_instance588();
    reg_declaration589 reg_declaration_instance589();
    reg_declaration590 reg_declaration_instance590();
    reg_declaration591 reg_declaration_instance591();
    reg_declaration592 reg_declaration_instance592();
    reg_declaration593 reg_declaration_instance593();
    reg_declaration594 reg_declaration_instance594();
    reg_declaration595 reg_declaration_instance595();
    reg_declaration596 reg_declaration_instance596();
    reg_declaration597 reg_declaration_instance597();
    reg_declaration598 reg_declaration_instance598();
    reg_declaration599 reg_declaration_instance599();
    reg_declaration600 reg_declaration_instance600();
    reg_declaration601 reg_declaration_instance601();
    reg_declaration602 reg_declaration_instance602();
    reg_declaration603 reg_declaration_instance603();
    reg_declaration604 reg_declaration_instance604();
    reg_declaration605 reg_declaration_instance605();
    reg_declaration606 reg_declaration_instance606();
    reg_declaration607 reg_declaration_instance607();
    reg_declaration608 reg_declaration_instance608();
    reg_declaration609 reg_declaration_instance609();
    reg_declaration610 reg_declaration_instance610();
    reg_declaration611 reg_declaration_instance611();
    reg_declaration612 reg_declaration_instance612();
    reg_declaration613 reg_declaration_instance613();
    reg_declaration614 reg_declaration_instance614();
    reg_declaration615 reg_declaration_instance615();
    reg_declaration616 reg_declaration_instance616();
    reg_declaration617 reg_declaration_instance617();
    reg_declaration618 reg_declaration_instance618();
    reg_declaration619 reg_declaration_instance619();
endmodule
//@
//author : andreib
module reg_declaration0;
reg abcd;
endmodule
//author : andreib
module reg_declaration1;
reg abcd , ABCD;
endmodule
//author : andreib
module reg_declaration2;
reg abcd , ABCD , _123;
endmodule
//author : andreib
module reg_declaration3;
reg abcd , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration4;
reg abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration5;
reg abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration6;
reg abcd , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration7;
reg abcd , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration8;
reg abcd , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration9;
reg abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration10;
reg abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration11;
reg abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration12;
reg abcd , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration13;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration14;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration15;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration16;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration17;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration18;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration19;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration20;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration21;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration22;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration23;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration24;
reg abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration25;
reg abcd , ABCD = 2;
endmodule
//author : andreib
module reg_declaration26;
reg abcd , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration27;
reg abcd , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration28;
reg abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration29;
reg abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration30;
reg abcd , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration31;
reg abcd [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration32;
reg abcd [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration33;
reg abcd [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration34;
reg abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration35;
reg abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration36;
reg abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration37;
reg abcd [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration38;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration39;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration40;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration41;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration42;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration43;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration44;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration45;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration46;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration47;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration48;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration49;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration50;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration51;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration52;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration53;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration54;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration55;
reg abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration56;
reg abcd [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration57;
reg abcd [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration58;
reg abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration59;
reg abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration60;
reg abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration61;
reg abcd [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration62;
reg abcd [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration63;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration64;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration65;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration66;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration67;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration68;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration69;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration70;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration71;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration72;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration73;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration74;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration75;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration76;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration77;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration78;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration79;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration80;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration81;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration82;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration83;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration84;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration85;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration86;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration87;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration88;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration89;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration90;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration91;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration92;
reg abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration93;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration94;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration95;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration96;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration97;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration98;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration99;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration100;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration101;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration102;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration103;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration104;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration105;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration106;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration107;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration108;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration109;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration110;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration111;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration112;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration113;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration114;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration115;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration116;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration117;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration118;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration119;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration120;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration121;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration122;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration123;
reg abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration124;
reg abcd = 2;
endmodule
//author : andreib
module reg_declaration125;
reg abcd = 2 , ABCD;
endmodule
//author : andreib
module reg_declaration126;
reg abcd = 2 , ABCD , _123;
endmodule
//author : andreib
module reg_declaration127;
reg abcd = 2 , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration128;
reg abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration129;
reg abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration130;
reg abcd = 2 , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration131;
reg abcd = 2 , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration132;
reg abcd = 2 , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration133;
reg abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration134;
reg abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration135;
reg abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration136;
reg abcd = 2 , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration137;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration138;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration139;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration140;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration141;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration142;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration143;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration144;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration145;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration146;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration147;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration148;
reg abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration149;
reg abcd = 2 , ABCD = 2;
endmodule
//author : andreib
module reg_declaration150;
reg abcd = 2 , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration151;
reg abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration152;
reg abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration153;
reg abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration154;
reg abcd = 2 , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration155;
reg [ 7 : 0 ] abcd;
endmodule
//author : andreib
module reg_declaration156;
reg [ 7 : 0 ] abcd , ABCD;
endmodule
//author : andreib
module reg_declaration157;
reg [ 7 : 0 ] abcd , ABCD , _123;
endmodule
//author : andreib
module reg_declaration158;
reg [ 7 : 0 ] abcd , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration159;
reg [ 7 : 0 ] abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration160;
reg [ 7 : 0 ] abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration161;
reg [ 7 : 0 ] abcd , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration162;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration163;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration164;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration165;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration166;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration167;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration168;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration169;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration170;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration171;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration172;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration173;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration174;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration175;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration176;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration177;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration178;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration179;
reg [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration180;
reg [ 7 : 0 ] abcd , ABCD = 2;
endmodule
//author : andreib
module reg_declaration181;
reg [ 7 : 0 ] abcd , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration182;
reg [ 7 : 0 ] abcd , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration183;
reg [ 7 : 0 ] abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration184;
reg [ 7 : 0 ] abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration185;
reg [ 7 : 0 ] abcd , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration186;
reg [ 7 : 0 ] abcd [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration187;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration188;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration189;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration190;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration191;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration192;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration193;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration194;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration195;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration196;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration197;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration198;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration199;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration200;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration201;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration202;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration203;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration204;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration205;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration206;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration207;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration208;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration209;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration210;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration211;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration212;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration213;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration214;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration215;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration216;
reg [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration217;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration218;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration219;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration220;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration221;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration222;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration223;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration224;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration225;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration226;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration227;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration228;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration229;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration230;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration231;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration232;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration233;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration234;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration235;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration236;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration237;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration238;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration239;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration240;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration241;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration242;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration243;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration244;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration245;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration246;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration247;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration248;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration249;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration250;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration251;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration252;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration253;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration254;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration255;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration256;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration257;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration258;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration259;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration260;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration261;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration262;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration263;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration264;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration265;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration266;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration267;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration268;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration269;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration270;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration271;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration272;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration273;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration274;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration275;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration276;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration277;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration278;
reg [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration279;
reg [ 7 : 0 ] abcd = 2;
endmodule
//author : andreib
module reg_declaration280;
reg [ 7 : 0 ] abcd = 2 , ABCD;
endmodule
//author : andreib
module reg_declaration281;
reg [ 7 : 0 ] abcd = 2 , ABCD , _123;
endmodule
//author : andreib
module reg_declaration282;
reg [ 7 : 0 ] abcd = 2 , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration283;
reg [ 7 : 0 ] abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration284;
reg [ 7 : 0 ] abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration285;
reg [ 7 : 0 ] abcd = 2 , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration286;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration287;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration288;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration289;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration290;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration291;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration292;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration293;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration294;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration295;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration296;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration297;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration298;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration299;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration300;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration301;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration302;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration303;
reg [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration304;
reg [ 7 : 0 ] abcd = 2 , ABCD = 2;
endmodule
//author : andreib
module reg_declaration305;
reg [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration306;
reg [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration307;
reg [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration308;
reg [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration309;
reg [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration310;
reg signed abcd;
endmodule
//author : andreib
module reg_declaration311;
reg signed abcd , ABCD;
endmodule
//author : andreib
module reg_declaration312;
reg signed abcd , ABCD , _123;
endmodule
//author : andreib
module reg_declaration313;
reg signed abcd , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration314;
reg signed abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration315;
reg signed abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration316;
reg signed abcd , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration317;
reg signed abcd , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration318;
reg signed abcd , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration319;
reg signed abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration320;
reg signed abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration321;
reg signed abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration322;
reg signed abcd , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration323;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration324;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration325;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration326;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration327;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration328;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration329;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration330;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration331;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration332;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration333;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration334;
reg signed abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration335;
reg signed abcd , ABCD = 2;
endmodule
//author : andreib
module reg_declaration336;
reg signed abcd , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration337;
reg signed abcd , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration338;
reg signed abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration339;
reg signed abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration340;
reg signed abcd , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration341;
reg signed abcd [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration342;
reg signed abcd [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration343;
reg signed abcd [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration344;
reg signed abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration345;
reg signed abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration346;
reg signed abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration347;
reg signed abcd [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration348;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration349;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration350;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration351;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration352;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration353;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration354;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration355;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration356;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration357;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration358;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration359;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration360;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration361;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration362;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration363;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration364;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration365;
reg signed abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration366;
reg signed abcd [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration367;
reg signed abcd [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration368;
reg signed abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration369;
reg signed abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration370;
reg signed abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration371;
reg signed abcd [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration372;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration373;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration374;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration375;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration376;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration377;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration378;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration379;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration380;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration381;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration382;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration383;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration384;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration385;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration386;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration387;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration388;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration389;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration390;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration391;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration392;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration393;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration394;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration395;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration396;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration397;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration398;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration399;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration400;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration401;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration402;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration403;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration404;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration405;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration406;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration407;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration408;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration409;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration410;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration411;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration412;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration413;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration414;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration415;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration416;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration417;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration418;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration419;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration420;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration421;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration422;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration423;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration424;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration425;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration426;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration427;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration428;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration429;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration430;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration431;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration432;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration433;
reg signed abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration434;
reg signed abcd = 2;
endmodule
//author : andreib
module reg_declaration435;
reg signed abcd = 2 , ABCD;
endmodule
//author : andreib
module reg_declaration436;
reg signed abcd = 2 , ABCD , _123;
endmodule
//author : andreib
module reg_declaration437;
reg signed abcd = 2 , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration438;
reg signed abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration439;
reg signed abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration440;
reg signed abcd = 2 , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration441;
reg signed abcd = 2 , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration442;
reg signed abcd = 2 , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration443;
reg signed abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration444;
reg signed abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration445;
reg signed abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration446;
reg signed abcd = 2 , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration447;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration448;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration449;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration450;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration451;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration452;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration453;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration454;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration455;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration456;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration457;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration458;
reg signed abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration459;
reg signed abcd = 2 , ABCD = 2;
endmodule
//author : andreib
module reg_declaration460;
reg signed abcd = 2 , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration461;
reg signed abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration462;
reg signed abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration463;
reg signed abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration464;
reg signed abcd = 2 , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration465;
reg signed [ 7 : 0 ] abcd;
endmodule
//author : andreib
module reg_declaration466;
reg signed [ 7 : 0 ] abcd , ABCD;
endmodule
//author : andreib
module reg_declaration467;
reg signed [ 7 : 0 ] abcd , ABCD , _123;
endmodule
//author : andreib
module reg_declaration468;
reg signed [ 7 : 0 ] abcd , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration469;
reg signed [ 7 : 0 ] abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration470;
reg signed [ 7 : 0 ] abcd , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration471;
reg signed [ 7 : 0 ] abcd , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration472;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration473;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration474;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration475;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration476;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration477;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration478;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration479;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration480;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration481;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration482;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration483;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration484;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration485;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration486;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration487;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration488;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration489;
reg signed [ 7 : 0 ] abcd , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration490;
reg signed [ 7 : 0 ] abcd , ABCD = 2;
endmodule
//author : andreib
module reg_declaration491;
reg signed [ 7 : 0 ] abcd , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration492;
reg signed [ 7 : 0 ] abcd , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration493;
reg signed [ 7 : 0 ] abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration494;
reg signed [ 7 : 0 ] abcd , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration495;
reg signed [ 7 : 0 ] abcd , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration496;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration497;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration498;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration499;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration500;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration501;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration502;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration503;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration504;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration505;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration506;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration507;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration508;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration509;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration510;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration511;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration512;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration513;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration514;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration515;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration516;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration517;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration518;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration519;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration520;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration521;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration522;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration523;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration524;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration525;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration526;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration527;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration528;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration529;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration530;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration531;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration532;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration533;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration534;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration535;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration536;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration537;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration538;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration539;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration540;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration541;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration542;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration543;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration544;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration545;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration546;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration547;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration548;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration549;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration550;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration551;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration552;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration553;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration554;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration555;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration556;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration557;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration558;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration559;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD;
endmodule
//author : andreib
module reg_declaration560;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123;
endmodule
//author : andreib
module reg_declaration561;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration562;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration563;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration564;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration565;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration566;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration567;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration568;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration569;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration570;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration571;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration572;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration573;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration574;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration575;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration576;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration577;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration578;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration579;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration580;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration581;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration582;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration583;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2;
endmodule
//author : andreib
module reg_declaration584;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration585;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration586;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration587;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration588;
reg signed [ 7 : 0 ] abcd [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , ABCD = 2 , _123 = 2;
endmodule
//author : andreib
module reg_declaration589;
reg signed [ 7 : 0 ] abcd = 2;
endmodule
//author : andreib
module reg_declaration590;
reg signed [ 7 : 0 ] abcd = 2 , ABCD;
endmodule
//author : andreib
module reg_declaration591;
reg signed [ 7 : 0 ] abcd = 2 , ABCD , _123;
endmodule
//author : andreib
module reg_declaration592;
reg signed [ 7 : 0 ] abcd = 2 , ABCD , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration593;
reg signed [ 7 : 0 ] abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration594;
reg signed [ 7 : 0 ] abcd = 2 , ABCD , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration595;
reg signed [ 7 : 0 ] abcd = 2 , ABCD , _123 = 2;
endmodule
//author : andreib
module reg_declaration596;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration597;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration598;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration599;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration600;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration601;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration602;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration603;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration604;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration605;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration606;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration607;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration608;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration609;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123;
endmodule
//author : andreib
module reg_declaration610;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration611;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration612;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration613;
reg signed [ 7 : 0 ] abcd = 2 , ABCD [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ] , _123 = 2;
endmodule
//author : andreib
module reg_declaration614;
reg signed [ 7 : 0 ] abcd = 2 , ABCD = 2;
endmodule
//author : andreib
module reg_declaration615;
reg signed [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123;
endmodule
//author : andreib
module reg_declaration616;
reg signed [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration617;
reg signed [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration618;
reg signed [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 [ 2 : 2 ] [ 2 : 2 ] [ 2 : 2 ];
endmodule
//author : andreib
module reg_declaration619;
reg signed [ 7 : 0 ] abcd = 2 , ABCD = 2 , _123 = 2;
endmodule
