-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u2_cslc_generated/code/vhdl/u2.vhd
-- FILE GENERATED ON : Mon Aug 31 07:19:47 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u2\ is
begin
end entity;

architecture \u2_logic\ of \u2\ is
  signal \x\ : csl_bit_vector(10#4# - 10#1# downto 10#0#);
  signal \clk\ : csl_bit;

  component \u1\ is
    port(\x\ : out csl_bit_vector(10#4# - 10#1# downto 10#0#);
         \clk\ : in csl_bit);
  end component;
begin
  -- In file 'TO BE IMPLEMENTED':14 instance name must difer from the instantiated obejct name.
end architecture;

