`include "defines.v"

module u4();
// Location of source csl unit: file name = ar16.csl line number = 47
  `include "u4.logic.v"
endmodule

