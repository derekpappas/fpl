// Test type: Decimal Numbers - z digit with underscore
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'dz__;
endmodule
