// Test type: Real numbers - exponent lower case sign
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=12.3e-12;
endmodule
