// Test type: Real numbers - real number with underscore
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=274.3_2_;
endmodule
