--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : z0.vh
--FILE GENERATED ON : Fri Aug 27 02:46:55 2010

a0.vhd
b0.vhd
c0.vhd
d0.vhd
e0.vhd
f0.vhd
g0.vhd
h0.vhd
i0.vhd
j0.vhd
k0.vhd
l0.vhd
m0.vhd
n0.vhd
o0.vhd
p0.vhd
q0.vhd
r0.vhd
s0.vhd
t0.vhd
u0.vhd
v0.vhd
w0.vhd
x0.vhd
y0.vhd
a1.vhd
b1.vhd
c1.vhd
d1.vhd
e1.vhd
f1.vhd
g1.vhd
h1.vhd
i1.vhd
j1.vhd
k1.vhd
l1.vhd
m1.vhd
n1.vhd
o1.vhd
p1.vhd
q1.vhd
r1.vhd
s1.vhd
t1.vhd
u1.vhd
v1.vhd
w1.vhd
x1.vhd
y1.vhd
z0.vhd
