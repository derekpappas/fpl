// Test type: seq_block - begin - block.id (ASCII) - 1 block item declaration - end
// Vparser rule name:
// Author: andreib
module seq_block7;
initial begin:abcdefghijklmnopqrstuvwxyzABCDEFGHIJKLMNOPQRSTUVWXYZ1234567890_$
	reg a;
	end
endmodule
