`include "Neuron_inc.v"

module Neuron_DW01_inc_8_0 ( A, SUM );
input  [7:0] A;
output [7:0] SUM;
    wire \carry[4] , \carry[2] , \carry[6] , \carry[7] , \carry[3] , 
        \carry[5] , n1;
    tri \A[7] , \A[6] , \A[4] , \A[0] , \A[3] , \A[2] , \A[5] , \A[1] ;
    assign \A[7]  = A[7];
    assign \A[6]  = A[6];
    assign \A[5]  = A[5];
    assign \A[4]  = A[4];
    assign \A[3]  = A[3];
    assign \A[2]  = A[2];
    assign \A[1]  = A[1];
    assign \A[0]  = A[0];
    GTECH_ADD_AB U1_1_3 ( .A(\A[3] ), .B(\carry[3] ), .S(SUM[3]), .COUT(
        \carry[4] ) );
    GTECH_ADD_AB U1_1_4 ( .A(\A[4] ), .B(\carry[4] ), .S(SUM[4]), .COUT(
        \carry[5] ) );
    GTECH_ADD_AB U1_1_1 ( .A(\A[1] ), .B(\A[0] ), .S(SUM[1]), .COUT(\carry[2] 
        ) );
    GTECH_ADD_AB U1_1_2 ( .A(\A[2] ), .B(\carry[2] ), .S(SUM[2]), .COUT(
        \carry[3] ) );
    GTECH_ADD_AB U1_1_5 ( .A(\A[5] ), .B(\carry[5] ), .S(SUM[5]), .COUT(
        \carry[6] ) );
    GTECH_ADD_AB U1_1_6 ( .A(\A[6] ), .B(\carry[6] ), .S(SUM[6]), .COUT(
        \carry[7] ) );
    GTECH_NOT U5 ( .A(\A[0] ), .Z(SUM[0]) );
    GTECH_OAI2N2 U6 ( .A(n1), .B(\A[7] ), .C(n1), .D(\A[7] ), .Z(SUM[7]) );
    GTECH_NOT U7 ( .A(\carry[7] ), .Z(n1) );
endmodule


module Neuron_DW02_mult_4_4_0 ( A, B, TC, PRODUCT );
input  [3:0] A;
input  [3:0] B;
output [7:0] PRODUCT;
input  TC;
    wire \CARRYB[2][1] , \ab[2][2] , \ab[2][0] , \ab[3][1] , \CARRYB[3][0] , 
        \ab[1][3] , \SUMB[1][2] , \ab[1][1] , \ab[0][2] , \SUMB[3][0] , 
        \CLA_CARRY[4] , \CARRYB[1][2] , \SUMB[3][2] , \SUMB[2][1] , 
        \CARRYB[1][0] , \CLA_SUM[5] , \ab[1][0] , \ab[0][3] , \CLA_SUM[4] , 
        \ab[1][2] , \CLA_CARRY[3] , \CARRYB[1][1] , \SUMB[3][1] , \SUMB[2][2] , 
        \ab[0][1] , \CARRYB[3][1] , \ab[3][2] , \ab[3][0] , \ab[2][3] , 
        \CARRYB[2][2] , \ab[2][1] , \SUMB[1][1] , \CARRYB[2][0] , n10, n11, 
        n12, n13, n14, n15, n16;
    GTECH_ADD_ABC S5_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\ab[2][3] ), 
        .S(\SUMB[3][2] ) );
    GTECH_ADD_ABC S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .C(\SUMB[1][2] 
        ), .S(\SUMB[2][1] ), .COUT(\CARRYB[2][1] ) );
    GTECH_ADD_ABC S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .C(\SUMB[1][1] 
        ), .S(PRODUCT[2]), .COUT(\CARRYB[2][0] ) );
    GTECH_ADD_ABC S4_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), 
        .S(\SUMB[3][1] ), .COUT(\CARRYB[3][1] ) );
    GTECH_ADD_ABC S14_3_2 ( .A(A[3]), .B(B[3]), .C(\SUMB[3][0] ), .S(PRODUCT
        [3]), .COUT(\CLA_CARRY[3] ) );
    GTECH_ADD_ABC S3_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .C(\ab[1][3] ), 
        .S(\SUMB[2][2] ), .COUT(\CARRYB[2][2] ) );
    GTECH_ADD_ABC S4_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), 
        .S(\SUMB[3][0] ), .COUT(\CARRYB[3][0] ) );
    GTECH_NOT U5 ( .A(n14), .Z(n16) );
    GTECH_AND_NOT U6 ( .A(\CARRYB[3][0] ), .B(n10), .Z(\CLA_CARRY[4] ) );
    GTECH_OAI2N2 U7 ( .A(\CARRYB[3][0] ), .B(n10), .C(\CARRYB[3][0] ), .D(n10), 
        .Z(\CLA_SUM[4] ) );
    GTECH_NOT U8 ( .A(\SUMB[3][1] ), .Z(n10) );
    GTECH_AND2 U9 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(\CARRYB[1][0] ) );
    GTECH_OAI2N2 U10 ( .A(n11), .B(\SUMB[3][2] ), .C(n11), .D(\SUMB[3][2] ), 
        .Z(\CLA_SUM[5] ) );
    GTECH_NOT U11 ( .A(\CARRYB[3][1] ), .Z(n11) );
    GTECH_AND_NOT U12 ( .A(\ab[1][2] ), .B(n12), .Z(\CARRYB[1][2] ) );
    GTECH_OAI2N2 U13 ( .A(\ab[1][2] ), .B(n12), .C(\ab[1][2] ), .D(n12), .Z(
        \SUMB[1][2] ) );
    GTECH_NOT U14 ( .A(\ab[0][3] ), .Z(n12) );
    GTECH_AND_NOT U15 ( .A(\ab[1][1] ), .B(n13), .Z(\CARRYB[1][1] ) );
    GTECH_OAI2N2 U16 ( .A(\ab[1][1] ), .B(n13), .C(\ab[1][1] ), .D(n13), .Z(
        \SUMB[1][1] ) );
    GTECH_NOT U17 ( .A(\ab[0][2] ), .Z(n13) );
    GTECH_AND_NOT U18 ( .A(A[3]), .B(B[2]), .Z(\ab[3][2] ) );
    GTECH_AND_NOT U19 ( .A(A[3]), .B(B[1]), .Z(\ab[3][1] ) );
    GTECH_AND_NOT U20 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
    GTECH_AND_NOT U21 ( .A(B[3]), .B(A[2]), .Z(\ab[2][3] ) );
    GTECH_AND2 U22 ( .A(A[2]), .B(B[2]), .Z(\ab[2][2] ) );
    GTECH_AND2 U23 ( .A(B[1]), .B(A[2]), .Z(\ab[2][1] ) );
    GTECH_AND2 U24 ( .A(B[0]), .B(A[2]), .Z(\ab[2][0] ) );
    GTECH_AND_NOT U25 ( .A(B[3]), .B(A[1]), .Z(\ab[1][3] ) );
    GTECH_AND2 U26 ( .A(A[1]), .B(B[2]), .Z(\ab[1][2] ) );
    GTECH_AND2 U27 ( .A(A[1]), .B(B[1]), .Z(\ab[1][1] ) );
    GTECH_AND2 U28 ( .A(B[0]), .B(A[1]), .Z(\ab[1][0] ) );
    GTECH_AND_NOT U29 ( .A(B[3]), .B(A[0]), .Z(\ab[0][3] ) );
    GTECH_AND2 U30 ( .A(B[2]), .B(A[0]), .Z(\ab[0][2] ) );
    GTECH_AND2 U31 ( .A(A[0]), .B(B[1]), .Z(\ab[0][1] ) );
    GTECH_AND_NOT U32 ( .A(n14), .B(n15), .Z(PRODUCT[4]) );
    GTECH_XOR3 U33 ( .A(\CLA_SUM[5] ), .B(\CLA_CARRY[4] ), .C(n16), .Z(PRODUCT
        [5]) );
    GTECH_NOR2 U34 ( .A(\CLA_SUM[4] ), .B(\CLA_CARRY[3] ), .Z(n15) );
    GTECH_NAND2 U35 ( .A(\CLA_SUM[4] ), .B(\CLA_CARRY[3] ), .Z(n14) );
endmodule


module Neuron ( .Variables({\Variables[0][-8][3] , \Variables[0][-8][2] , 
    \Variables[0][-8][1] , \Variables[0][-8][0] , \Variables[0][-7][3] , 
    \Variables[0][-7][2] , \Variables[0][-7][1] , \Variables[0][-7][0] , 
    \Variables[0][-6][3] , \Variables[0][-6][2] , \Variables[0][-6][1] , 
    \Variables[0][-6][0] , \Variables[0][-5][3] , \Variables[0][-5][2] , 
    \Variables[0][-5][1] , \Variables[0][-5][0] , \Variables[0][-4][3] , 
    \Variables[0][-4][2] , \Variables[0][-4][1] , \Variables[0][-4][0] , 
    \Variables[0][-3][3] , \Variables[0][-3][2] , \Variables[0][-3][1] , 
    \Variables[0][-3][0] , \Variables[0][-2][3] , \Variables[0][-2][2] , 
    \Variables[0][-2][1] , \Variables[0][-2][0] , \Variables[0][-1][3] , 
    \Variables[0][-1][2] , \Variables[0][-1][1] , \Variables[0][-1][0] , 
    \Variables[0][0][3] , \Variables[0][0][2] , \Variables[0][0][1] , 
    \Variables[0][0][0] , \Variables[0][1][3] , \Variables[0][1][2] , 
    \Variables[0][1][1] , \Variables[0][1][0] , \Variables[0][2][3] , 
    \Variables[0][2][2] , \Variables[0][2][1] , \Variables[0][2][0] , 
    \Variables[0][3][3] , \Variables[0][3][2] , \Variables[0][3][1] , 
    \Variables[0][3][0] , \Variables[0][4][3] , \Variables[0][4][2] , 
    \Variables[0][4][1] , \Variables[0][4][0] , \Variables[0][5][3] , 
    \Variables[0][5][2] , \Variables[0][5][1] , \Variables[0][5][0] , 
    \Variables[0][6][3] , \Variables[0][6][2] , \Variables[0][6][1] , 
    \Variables[0][6][0] , \Variables[0][7][3] , \Variables[0][7][2] , 
    \Variables[0][7][1] , \Variables[0][7][0] , \Variables[1][-8][3] , 
    \Variables[1][-8][2] , \Variables[1][-8][1] , \Variables[1][-8][0] , 
    \Variables[1][-7][3] , \Variables[1][-7][2] , \Variables[1][-7][1] , 
    \Variables[1][-7][0] , \Variables[1][-6][3] , \Variables[1][-6][2] , 
    \Variables[1][-6][1] , \Variables[1][-6][0] , \Variables[1][-5][3] , 
    \Variables[1][-5][2] , \Variables[1][-5][1] , \Variables[1][-5][0] , 
    \Variables[1][-4][3] , \Variables[1][-4][2] , \Variables[1][-4][1] , 
    \Variables[1][-4][0] , \Variables[1][-3][3] , \Variables[1][-3][2] , 
    \Variables[1][-3][1] , \Variables[1][-3][0] , \Variables[1][-2][3] , 
    \Variables[1][-2][2] , \Variables[1][-2][1] , \Variables[1][-2][0] , 
    \Variables[1][-1][3] , \Variables[1][-1][2] , \Variables[1][-1][1] , 
    \Variables[1][-1][0] , \Variables[1][0][3] , \Variables[1][0][2] , 
    \Variables[1][0][1] , \Variables[1][0][0] , \Variables[1][1][3] , 
    \Variables[1][1][2] , \Variables[1][1][1] , \Variables[1][1][0] , 
    \Variables[1][2][3] , \Variables[1][2][2] , \Variables[1][2][1] , 
    \Variables[1][2][0] , \Variables[1][3][3] , \Variables[1][3][2] , 
    \Variables[1][3][1] , \Variables[1][3][0] , \Variables[1][4][3] , 
    \Variables[1][4][2] , \Variables[1][4][1] , \Variables[1][4][0] , 
    \Variables[1][5][3] , \Variables[1][5][2] , \Variables[1][5][1] , 
    \Variables[1][5][0] , \Variables[1][6][3] , \Variables[1][6][2] , 
    \Variables[1][6][1] , \Variables[1][6][0] , \Variables[1][7][3] , 
    \Variables[1][7][2] , \Variables[1][7][1] , \Variables[1][7][0] , 
    \Variables[2][-8][3] , \Variables[2][-8][2] , \Variables[2][-8][1] , 
    \Variables[2][-8][0] , \Variables[2][-7][3] , \Variables[2][-7][2] , 
    \Variables[2][-7][1] , \Variables[2][-7][0] , \Variables[2][-6][3] , 
    \Variables[2][-6][2] , \Variables[2][-6][1] , \Variables[2][-6][0] , 
    \Variables[2][-5][3] , \Variables[2][-5][2] , \Variables[2][-5][1] , 
    \Variables[2][-5][0] , \Variables[2][-4][3] , \Variables[2][-4][2] , 
    \Variables[2][-4][1] , \Variables[2][-4][0] , \Variables[2][-3][3] , 
    \Variables[2][-3][2] , \Variables[2][-3][1] , \Variables[2][-3][0] , 
    \Variables[2][-2][3] , \Variables[2][-2][2] , \Variables[2][-2][1] , 
    \Variables[2][-2][0] , \Variables[2][-1][3] , \Variables[2][-1][2] , 
    \Variables[2][-1][1] , \Variables[2][-1][0] , \Variables[2][0][3] , 
    \Variables[2][0][2] , \Variables[2][0][1] , \Variables[2][0][0] , 
    \Variables[2][1][3] , \Variables[2][1][2] , \Variables[2][1][1] , 
    \Variables[2][1][0] , \Variables[2][2][3] , \Variables[2][2][2] , 
    \Variables[2][2][1] , \Variables[2][2][0] , \Variables[2][3][3] , 
    \Variables[2][3][2] , \Variables[2][3][1] , \Variables[2][3][0] , 
    \Variables[2][4][3] , \Variables[2][4][2] , \Variables[2][4][1] , 
    \Variables[2][4][0] , \Variables[2][5][3] , \Variables[2][5][2] , 
    \Variables[2][5][1] , \Variables[2][5][0] , \Variables[2][6][3] , 
    \Variables[2][6][2] , \Variables[2][6][1] , \Variables[2][6][0] , 
    \Variables[2][7][3] , \Variables[2][7][2] , \Variables[2][7][1] , 
    \Variables[2][7][0] , \Variables[3][-8][3] , \Variables[3][-8][2] , 
    \Variables[3][-8][1] , \Variables[3][-8][0] , \Variables[3][-7][3] , 
    \Variables[3][-7][2] , \Variables[3][-7][1] , \Variables[3][-7][0] , 
    \Variables[3][-6][3] , \Variables[3][-6][2] , \Variables[3][-6][1] , 
    \Variables[3][-6][0] , \Variables[3][-5][3] , \Variables[3][-5][2] , 
    \Variables[3][-5][1] , \Variables[3][-5][0] , \Variables[3][-4][3] , 
    \Variables[3][-4][2] , \Variables[3][-4][1] , \Variables[3][-4][0] , 
    \Variables[3][-3][3] , \Variables[3][-3][2] , \Variables[3][-3][1] , 
    \Variables[3][-3][0] , \Variables[3][-2][3] , \Variables[3][-2][2] , 
    \Variables[3][-2][1] , \Variables[3][-2][0] , \Variables[3][-1][3] , 
    \Variables[3][-1][2] , \Variables[3][-1][1] , \Variables[3][-1][0] , 
    \Variables[3][0][3] , \Variables[3][0][2] , \Variables[3][0][1] , 
    \Variables[3][0][0] , \Variables[3][1][3] , \Variables[3][1][2] , 
    \Variables[3][1][1] , \Variables[3][1][0] , \Variables[3][2][3] , 
    \Variables[3][2][2] , \Variables[3][2][1] , \Variables[3][2][0] , 
    \Variables[3][3][3] , \Variables[3][3][2] , \Variables[3][3][1] , 
    \Variables[3][3][0] , \Variables[3][4][3] , \Variables[3][4][2] , 
    \Variables[3][4][1] , \Variables[3][4][0] , \Variables[3][5][3] , 
    \Variables[3][5][2] , \Variables[3][5][1] , \Variables[3][5][0] , 
    \Variables[3][6][3] , \Variables[3][6][2] , \Variables[3][6][1] , 
    \Variables[3][6][0] , \Variables[3][7][3] , \Variables[3][7][2] , 
    \Variables[3][7][1] , \Variables[3][7][0] , \Variables[4][-8][3] , 
    \Variables[4][-8][2] , \Variables[4][-8][1] , \Variables[4][-8][0] , 
    \Variables[4][-7][3] , \Variables[4][-7][2] , \Variables[4][-7][1] , 
    \Variables[4][-7][0] , \Variables[4][-6][3] , \Variables[4][-6][2] , 
    \Variables[4][-6][1] , \Variables[4][-6][0] , \Variables[4][-5][3] , 
    \Variables[4][-5][2] , \Variables[4][-5][1] , \Variables[4][-5][0] , 
    \Variables[4][-4][3] , \Variables[4][-4][2] , \Variables[4][-4][1] , 
    \Variables[4][-4][0] , \Variables[4][-3][3] , \Variables[4][-3][2] , 
    \Variables[4][-3][1] , \Variables[4][-3][0] , \Variables[4][-2][3] , 
    \Variables[4][-2][2] , \Variables[4][-2][1] , \Variables[4][-2][0] , 
    \Variables[4][-1][3] , \Variables[4][-1][2] , \Variables[4][-1][1] , 
    \Variables[4][-1][0] , \Variables[4][0][3] , \Variables[4][0][2] , 
    \Variables[4][0][1] , \Variables[4][0][0] , \Variables[4][1][3] , 
    \Variables[4][1][2] , \Variables[4][1][1] , \Variables[4][1][0] , 
    \Variables[4][2][3] , \Variables[4][2][2] , \Variables[4][2][1] , 
    \Variables[4][2][0] , \Variables[4][3][3] , \Variables[4][3][2] , 
    \Variables[4][3][1] , \Variables[4][3][0] , \Variables[4][4][3] , 
    \Variables[4][4][2] , \Variables[4][4][1] , \Variables[4][4][0] , 
    \Variables[4][5][3] , \Variables[4][5][2] , \Variables[4][5][1] , 
    \Variables[4][5][0] , \Variables[4][6][3] , \Variables[4][6][2] , 
    \Variables[4][6][1] , \Variables[4][6][0] , \Variables[4][7][3] , 
    \Variables[4][7][2] , \Variables[4][7][1] , \Variables[4][7][0] }), 
    InstructionPtr, MemoryPtr, MemoryWriteValue, MemoryReadValue, Read, Write, 
    MemoryReady, .NextInstruction({\NextInstruction[INSTRUCTION][0] , 
    \NextInstruction[INSTRUCTION][1] , \NextInstruction[INSTRUCTION][2] , 
    \NextInstruction[INSTRUCTION][3] , \NextInstruction[PARAMETER][3] , 
    \NextInstruction[PARAMETER][2] , \NextInstruction[PARAMETER][1] , 
    \NextInstruction[PARAMETER][0] }), IRQ, InstructionReady, clk, Reset );
inout  [7:0] InstructionPtr;
inout  [7:0] MemoryPtr;
output [7:0] MemoryWriteValue;
input  [7:0] MemoryReadValue;
inout  [0:4] IRQ;
input  MemoryReady, \NextInstruction[INSTRUCTION][0] , 
    \NextInstruction[INSTRUCTION][1] , \NextInstruction[INSTRUCTION][2] , 
    \NextInstruction[INSTRUCTION][3] , \NextInstruction[PARAMETER][3] , 
    \NextInstruction[PARAMETER][2] , \NextInstruction[PARAMETER][1] , 
    \NextInstruction[PARAMETER][0] , InstructionReady, clk, Reset;
inout  \Variables[0][-8][3] , \Variables[0][-8][2] , \Variables[0][-8][1] , 
    \Variables[0][-8][0] , \Variables[0][-7][3] , \Variables[0][-7][2] , 
    \Variables[0][-7][1] , \Variables[0][-7][0] , \Variables[0][-6][3] , 
    \Variables[0][-6][2] , \Variables[0][-6][1] , \Variables[0][-6][0] , 
    \Variables[0][-5][3] , \Variables[0][-5][2] , \Variables[0][-5][1] , 
    \Variables[0][-5][0] , \Variables[0][-4][3] , \Variables[0][-4][2] , 
    \Variables[0][-4][1] , \Variables[0][-4][0] , \Variables[0][-3][3] , 
    \Variables[0][-3][2] , \Variables[0][-3][1] , \Variables[0][-3][0] , 
    \Variables[0][-2][3] , \Variables[0][-2][2] , \Variables[0][-2][1] , 
    \Variables[0][-2][0] , \Variables[0][-1][3] , \Variables[0][-1][2] , 
    \Variables[0][-1][1] , \Variables[0][-1][0] , \Variables[0][0][3] , 
    \Variables[0][0][2] , \Variables[0][0][1] , \Variables[0][0][0] , 
    \Variables[0][1][3] , \Variables[0][1][2] , \Variables[0][1][1] , 
    \Variables[0][1][0] , \Variables[0][2][3] , \Variables[0][2][2] , 
    \Variables[0][2][1] , \Variables[0][2][0] , \Variables[0][3][3] , 
    \Variables[0][3][2] , \Variables[0][3][1] , \Variables[0][3][0] , 
    \Variables[0][4][3] , \Variables[0][4][2] , \Variables[0][4][1] , 
    \Variables[0][4][0] , \Variables[0][5][3] , \Variables[0][5][2] , 
    \Variables[0][5][1] , \Variables[0][5][0] , \Variables[0][6][3] , 
    \Variables[0][6][2] , \Variables[0][6][1] , \Variables[0][6][0] , 
    \Variables[0][7][3] , \Variables[0][7][2] , \Variables[0][7][1] , 
    \Variables[0][7][0] , \Variables[1][-8][3] , \Variables[1][-8][2] , 
    \Variables[1][-8][1] , \Variables[1][-8][0] , \Variables[1][-7][3] , 
    \Variables[1][-7][2] , \Variables[1][-7][1] , \Variables[1][-7][0] , 
    \Variables[1][-6][3] , \Variables[1][-6][2] , \Variables[1][-6][1] , 
    \Variables[1][-6][0] , \Variables[1][-5][3] , \Variables[1][-5][2] , 
    \Variables[1][-5][1] , \Variables[1][-5][0] , \Variables[1][-4][3] , 
    \Variables[1][-4][2] , \Variables[1][-4][1] , \Variables[1][-4][0] , 
    \Variables[1][-3][3] , \Variables[1][-3][2] , \Variables[1][-3][1] , 
    \Variables[1][-3][0] , \Variables[1][-2][3] , \Variables[1][-2][2] , 
    \Variables[1][-2][1] , \Variables[1][-2][0] , \Variables[1][-1][3] , 
    \Variables[1][-1][2] , \Variables[1][-1][1] , \Variables[1][-1][0] , 
    \Variables[1][0][3] , \Variables[1][0][2] , \Variables[1][0][1] , 
    \Variables[1][0][0] , \Variables[1][1][3] , \Variables[1][1][2] , 
    \Variables[1][1][1] , \Variables[1][1][0] , \Variables[1][2][3] , 
    \Variables[1][2][2] , \Variables[1][2][1] , \Variables[1][2][0] , 
    \Variables[1][3][3] , \Variables[1][3][2] , \Variables[1][3][1] , 
    \Variables[1][3][0] , \Variables[1][4][3] , \Variables[1][4][2] , 
    \Variables[1][4][1] , \Variables[1][4][0] , \Variables[1][5][3] , 
    \Variables[1][5][2] , \Variables[1][5][1] , \Variables[1][5][0] , 
    \Variables[1][6][3] , \Variables[1][6][2] , \Variables[1][6][1] , 
    \Variables[1][6][0] , \Variables[1][7][3] , \Variables[1][7][2] , 
    \Variables[1][7][1] , \Variables[1][7][0] , \Variables[2][-8][3] , 
    \Variables[2][-8][2] , \Variables[2][-8][1] , \Variables[2][-8][0] , 
    \Variables[2][-7][3] , \Variables[2][-7][2] , \Variables[2][-7][1] , 
    \Variables[2][-7][0] , \Variables[2][-6][3] , \Variables[2][-6][2] , 
    \Variables[2][-6][1] , \Variables[2][-6][0] , \Variables[2][-5][3] , 
    \Variables[2][-5][2] , \Variables[2][-5][1] , \Variables[2][-5][0] , 
    \Variables[2][-4][3] , \Variables[2][-4][2] , \Variables[2][-4][1] , 
    \Variables[2][-4][0] , \Variables[2][-3][3] , \Variables[2][-3][2] , 
    \Variables[2][-3][1] , \Variables[2][-3][0] , \Variables[2][-2][3] , 
    \Variables[2][-2][2] , \Variables[2][-2][1] , \Variables[2][-2][0] , 
    \Variables[2][-1][3] , \Variables[2][-1][2] , \Variables[2][-1][1] , 
    \Variables[2][-1][0] , \Variables[2][0][3] , \Variables[2][0][2] , 
    \Variables[2][0][1] , \Variables[2][0][0] , \Variables[2][1][3] , 
    \Variables[2][1][2] , \Variables[2][1][1] , \Variables[2][1][0] , 
    \Variables[2][2][3] , \Variables[2][2][2] , \Variables[2][2][1] , 
    \Variables[2][2][0] , \Variables[2][3][3] , \Variables[2][3][2] , 
    \Variables[2][3][1] , \Variables[2][3][0] , \Variables[2][4][3] , 
    \Variables[2][4][2] , \Variables[2][4][1] , \Variables[2][4][0] , 
    \Variables[2][5][3] , \Variables[2][5][2] , \Variables[2][5][1] , 
    \Variables[2][5][0] , \Variables[2][6][3] , \Variables[2][6][2] , 
    \Variables[2][6][1] , \Variables[2][6][0] , \Variables[2][7][3] , 
    \Variables[2][7][2] , \Variables[2][7][1] , \Variables[2][7][0] , 
    \Variables[3][-8][3] , \Variables[3][-8][2] , \Variables[3][-8][1] , 
    \Variables[3][-8][0] , \Variables[3][-7][3] , \Variables[3][-7][2] , 
    \Variables[3][-7][1] , \Variables[3][-7][0] , \Variables[3][-6][3] , 
    \Variables[3][-6][2] , \Variables[3][-6][1] , \Variables[3][-6][0] , 
    \Variables[3][-5][3] , \Variables[3][-5][2] , \Variables[3][-5][1] , 
    \Variables[3][-5][0] , \Variables[3][-4][3] , \Variables[3][-4][2] , 
    \Variables[3][-4][1] , \Variables[3][-4][0] , \Variables[3][-3][3] , 
    \Variables[3][-3][2] , \Variables[3][-3][1] , \Variables[3][-3][0] , 
    \Variables[3][-2][3] , \Variables[3][-2][2] , \Variables[3][-2][1] , 
    \Variables[3][-2][0] , \Variables[3][-1][3] , \Variables[3][-1][2] , 
    \Variables[3][-1][1] , \Variables[3][-1][0] , \Variables[3][0][3] , 
    \Variables[3][0][2] , \Variables[3][0][1] , \Variables[3][0][0] , 
    \Variables[3][1][3] , \Variables[3][1][2] , \Variables[3][1][1] , 
    \Variables[3][1][0] , \Variables[3][2][3] , \Variables[3][2][2] , 
    \Variables[3][2][1] , \Variables[3][2][0] , \Variables[3][3][3] , 
    \Variables[3][3][2] , \Variables[3][3][1] , \Variables[3][3][0] , 
    \Variables[3][4][3] , \Variables[3][4][2] , \Variables[3][4][1] , 
    \Variables[3][4][0] , \Variables[3][5][3] , \Variables[3][5][2] , 
    \Variables[3][5][1] , \Variables[3][5][0] , \Variables[3][6][3] , 
    \Variables[3][6][2] , \Variables[3][6][1] , \Variables[3][6][0] , 
    \Variables[3][7][3] , \Variables[3][7][2] , \Variables[3][7][1] , 
    \Variables[3][7][0] , \Variables[4][-8][3] , \Variables[4][-8][2] , 
    \Variables[4][-8][1] , \Variables[4][-8][0] , \Variables[4][-7][3] , 
    \Variables[4][-7][2] , \Variables[4][-7][1] , \Variables[4][-7][0] , 
    \Variables[4][-6][3] , \Variables[4][-6][2] , \Variables[4][-6][1] , 
    \Variables[4][-6][0] , \Variables[4][-5][3] , \Variables[4][-5][2] , 
    \Variables[4][-5][1] , \Variables[4][-5][0] , \Variables[4][-4][3] , 
    \Variables[4][-4][2] , \Variables[4][-4][1] , \Variables[4][-4][0] , 
    \Variables[4][-3][3] , \Variables[4][-3][2] , \Variables[4][-3][1] , 
    \Variables[4][-3][0] , \Variables[4][-2][3] , \Variables[4][-2][2] , 
    \Variables[4][-2][1] , \Variables[4][-2][0] , \Variables[4][-1][3] , 
    \Variables[4][-1][2] , \Variables[4][-1][1] , \Variables[4][-1][0] , 
    \Variables[4][0][3] , \Variables[4][0][2] , \Variables[4][0][1] , 
    \Variables[4][0][0] , \Variables[4][1][3] , \Variables[4][1][2] , 
    \Variables[4][1][1] , \Variables[4][1][0] , \Variables[4][2][3] , 
    \Variables[4][2][2] , \Variables[4][2][1] , \Variables[4][2][0] , 
    \Variables[4][3][3] , \Variables[4][3][2] , \Variables[4][3][1] , 
    \Variables[4][3][0] , \Variables[4][4][3] , \Variables[4][4][2] , 
    \Variables[4][4][1] , \Variables[4][4][0] , \Variables[4][5][3] , 
    \Variables[4][5][2] , \Variables[4][5][1] , \Variables[4][5][0] , 
    \Variables[4][6][3] , \Variables[4][6][2] , \Variables[4][6][1] , 
    \Variables[4][6][0] , \Variables[4][7][3] , \Variables[4][7][2] , 
    \Variables[4][7][1] , \Variables[4][7][0] , Read, Write;
    wire \Variables2830[3][-7][3] , InterruptJump, \InstructionPtr3995[6] , 
        IRQWait611, \Variables2830[3][-3][1] , \ClockCycleCount621[1] , 
        \Answer2629[0] , n658, \Variables2830[0][-3][0] , 
        \Variables2830[1][1][2] , \Variables2830[3][2][3] , \sum1105[0] , 
        \Variables2830[0][-7][2] , \Variables2830[3][6][1] , n_693, 
        \Variables2830[1][5][0] , \Variables2830[4][-8][1] , 
        \Variables2830[3][-2][2] , ReturnJump, 
        \RegularWriteRegister_Index848[2] , \Variables2830[3][-6][0] , 
        \MemoryPtr3672[7] , \Answer639[1] , \Variables2830[0][-6][1] , 
        \Variables2830[1][4][3] , \Variables2830[3][7][2] , 
        \Variables2830[0][-2][3] , \Variables2830[3][3][0] , 
        \Variables2830[1][0][1] , \Variables2830[1][-1][1] , IRQCLKEnable676, 
        \Variables2830[1][-5][3] , OutOfRangeException2645, 
        \Variables2830[4][-6][1] , \Variables2830[4][0][0] , 
        \Variables2830[0][5][3] , \Variables2830[2][6][2] , Condition, 
        \Variables2830[2][-5][2] , \IPRELOAD_Index[2] , 
        \Variables2830[2][-1][0] , \Variables2830[2][2][0] , 
        \Variables2830[0][1][1] , \InstructionPtr3995[2] , \IRQ_Index[2] , 
        \Variables2830[4][-2][3] , \Variables2830[4][4][2] , 
        \Variables2830[1][-4][0] , \Variables2830[3][-8][0] , RegularJump, 
        ResetStarted, \Variables2830[4][5][1] , \Variables2830[4][-3][0] , 
        \MemoryPtr3672[3] , \Variables2830[0][0][2] , \Variables2830[2][3][3] , 
        n603, \Variables2830[2][-4][1] , \Variables2830[2][7][1] , 
        \Variables2830[0][-8][1] , \Variables2830[0][4][0] , 
        \Variables2830[4][-7][2] , \Variables2830[4][1][3] , 
        \Variables2830[4][-3][2] , \MemoryPtr3672[1] , 
        \Variables2830[4][5][3] , \Variables2830[2][3][1] , 
        \Variables2830[0][0][0] , \Variables2830[0][4][2] , 
        \Variables2830[0][-8][3] , \Variables2830[2][-4][3] , 
        \Variables2830[2][7][3] , \Variables2830[4][-7][0] , 
        \Variables2830[4][1][1] , \Variables2830[3][-8][2] , 
        \Variables2830[1][-4][2] , \Variables2830[4][-6][3] , 
        \Variables2830[4][0][2] , \Variables2830[2][-5][0] , 
        \Variables2830[2][6][0] , \Variables2830[0][5][1] , 
        \Variables2830[0][1][3] , \Variables2830[2][2][2] , 
        \Variables2830[2][-1][2] , \InstructionPtr3995[0] , 
        \Variables2830[4][-2][1] , \IRQ_Index[0] , \Variables2830[4][4][0] , 
        \Variables2830[1][-1][3] , \ClockCycleCount[1] , 
        \Variables2830[1][-5][1] , \Answer639[3] , \Variables2830[0][-6][3] , 
        RegularRegisterWrite, \Variables2830[3][7][0] , 
        \Variables2830[1][4][1] , \Variables2830[0][-2][1] , 
        \Variables2830[1][0][3] , \Variables2830[3][3][2] , IRQEnable685, n686, 
        \Variables2830[3][-2][0] , \n630[3] , 
        \RegularWriteRegister_Index848[0] , \n668[3] , 
        \Variables2830[3][-6][2] , \MemoryPtr3672[5] , 
        \Variables2830[0][-3][2] , \Variables2830[3][2][1] , 
        \Variables2830[1][1][0] , \sum1105[2] , \Variables2830[0][-7][0] , 
        \Variables2830[1][5][2] , \Variables2830[3][6][3] , 
        \Variables2830[4][-8][3] , \Variables2830[3][-7][1] , 
        \InstructionPtr3995[4] , n_566, \Variables2830[3][-3][3] , 
        \Answer2629[2] , n_452, \Variables2830[4][6][2] , \product1846[5] , 
        \IPRELOAD_Table[1] , n_358, \Variables2830[2][-3][0] , 
        \Variables2830[2][0][0] , \RegularWriteRegister_Index[3] , 
        \Variables2830[0][3][1] , \Variables2830[0][7][3] , 
        \Variables2830[2][-7][2] , \Variables2830[2][4][2] , 
        \Variables2830[4][2][0] , \Variables2830[4][-4][1] , 
        \CycleWaveform34[3] , \Variables2830[1][-7][3] , \TableSelect667[2] , 
        \Variables2830[1][-3][1] , \Variables2830[4][3][3] , 
        \Variables2830[4][-5][2] , \sum2964[3] , \Variables2830[2][5][1] , 
        \Variables2830[2][-6][1] , \Variables2830[0][6][0] , 
        \Variables2830[0][2][2] , \Variables2830[2][1][3] , 
        \Variables2830[2][-2][3] , \Variables2830[4][7][1] , 
        \Variables2830[4][-1][0] , n_168, \Variables2830[1][-2][2] , 
        \Variables2830[1][-6][0] , \n3996[7] , \Variables2830[3][4][1] , 
        \Variables2830[1][7][0] , \n706[3] , \Variables2830[0][-5][2] , 
        \Variables2830[1][3][2] , \Variables2830[3][0][3] , 
        \Variables2830[0][-1][0] , \Upper[2] , \Variables2830[3][-1][1] , 
        \IPRELOAD_Index3559[2] , \Variables2830[3][-5][3] , 
        \Variables2830[1][2][1] , \Variables2830[3][1][0] , \CycleWaveform[2] , 
        n_324, \Variables2830[1][6][3] , \Variables2830[3][5][2] , 
        \Variables2830[0][-4][1] , \Variables2830[2][-8][1] , IRQCLKEnable, 
        \Lower[1] , \Variables2830[3][-4][0] , \Variables2830[1][-8][0] , 
        \sum2964[7] , IRQInProcess602, \Lower[3] , \Variables2830[1][-8][2] , 
        \Variables2830[3][-4][2] , \sum2964[5] , n_689, 
        \Variables2830[1][2][3] , \Variables2830[3][1][2] , \IRQ2736[4] , 
        \Variables2830[3][5][0] , \Variables2830[1][6][1] , 
        \Exception_Index[3] , \Variables2830[2][-8][3] , 
        \IPRELOAD_Table3551[2] , \Variables2830[0][-4][3] , n_323, 
        \n2831[0][-8][3] , \Upper[0] , \Variables2830[3][-1][3] , 
        \IPRELOAD_Index3559[0] , n_692, \Variables2830[3][-5][1] , 
        \product1846[3] , \CycleWaveform[4] , \Variables2830[1][7][2] , 
        \Variables2830[3][4][3] , \Variables2830[0][-5][0] , 
        \Variables2830[1][3][0] , \Variables2830[3][0][1] , 
        \Variables2830[0][-1][2] , \CycleWaveform34[5] , 
        \Variables2830[1][-2][0] , \Variables2830[1][-6][2] , n3641, 
        \Variables2830[4][3][1] , \Variables2830[4][-5][0] , \sum2964[1] , 
        \Variables2830[0][6][2] , \Variables2830[2][5][3] , 
        \Variables2830[2][-6][3] , \Variables2830[2][-2][1] , 
        \Variables2830[2][1][1] , \Variables2830[0][2][0] , 
        \Variables2830[4][7][3] , \Variables2830[4][-1][2] , 
        \CycleWaveform34[1] , \Variables2830[1][-7][1] , n677, 
        \TableSelect667[0] , \CycleWaveform[5] , \Variables2830[1][-3][3] , 
        \Variables2830[4][6][0] , \Variables2830[0][3][3] , 
        \RegularWriteRegister_Index[1] , \Variables2830[2][-3][2] , 
        \Variables2830[2][0][2] , \TableSelect[0] , \Variables2830[2][-7][0] , 
        \Variables2830[2][4][0] , \Variables2830[0][7][1] , 
        \Variables2830[4][2][2] , \Variables2830[4][-4][3] , n612, 
        \Variables2830[1][-2][1] , \Variables2830[1][-6][3] , \sum2964[0] , 
        \Variables2830[2][-6][2] , \Variables2830[2][5][2] , 
        \Variables2830[0][6][3] , IRQInProcess, \Variables2830[4][3][0] , 
        n_690, \Variables2830[4][-5][1] , \Variables2830[4][7][2] , 
        \Variables2830[4][-1][3] , \Variables2830[0][2][1] , 
        \Variables2830[2][-2][0] , \Variables2830[2][1][0] , 
        \CycleWaveform34[0] , \Variables2830[1][-7][0] , 
        \Variables2830[1][-3][2] , \TableSelect667[1] , \CycleWaveform[1] , 
        \IPRELOAD_Table[2] , \Variables2830[0][3][2] , 
        \Variables2830[2][-3][3] , \Variables2830[2][0][3] , 
        \RegularWriteRegister_Index[0] , \Variables2830[4][6][1] , 
        \n2831[0][-3][3] , \Variables2830[4][2][3] , \Variables2830[4][-4][2] , 
        \TableSelect[1] , \Variables2830[0][7][0] , \Variables2830[2][4][1] , 
        \Variables2830[2][-7][1] , \Lower[2] , \Variables2830[3][-4][3] , 
        \Variables2830[1][-8][3] , IRQJump, \sum2964[4] , 
        \Variables2830[3][1][3] , \Variables2830[1][2][2] , 
        \Variables2830[1][6][0] , \Variables2830[3][5][1] , 
        \Variables2830[2][-8][2] , \Exception_Index[2] , 
        \Variables2830[0][-4][2] , \IPRELOAD_Index3559[1] , \Upper[1] , 
        \Variables2830[3][-1][2] , \product1846[2] , \Variables2830[3][-5][0] , 
        \n640[3] , \Variables2830[3][4][2] , \Variables2830[1][7][3] , 
        \Variables2830[0][-5][1] , \CycleWaveform34[4] , 
        \Variables2830[1][3][1] , \Variables2830[3][0][0] , 
        \Variables2830[0][-1][3] , \Variables2830[1][7][1] , 
        \Variables2830[3][4][0] , \Variables2830[0][-5][3] , \n3651[7] , n_660, 
        \Variables2830[3][0][2] , \Variables2830[1][3][3] , 
        \Variables2830[0][-1][1] , \IPRELOAD_Index3559[3] , \Upper[3] , 
        \CycleWaveform[3] , \Variables2830[3][-1][0] , 
        \Variables2830[3][-5][2] , \Variables2830[1][2][0] , 
        \Variables2830[3][1][1] , n_398, \Variables2830[3][5][3] , 
        \Variables2830[1][6][2] , \Variables2830[0][-4][0] , 
        \Variables2830[2][-8][0] , \Exception_Index[0] , 
        \IPRELOAD_Table3551[1] , \Lower[0] , \Variables2830[3][-4][1] , 
        \Variables2830[1][-8][1] , n_4166, \sum2964[6] , \IPRELOAD_Table[0] , 
        \RegularWriteRegister_Index[2] , \Variables2830[0][3][0] , 
        \Variables2830[2][-3][1] , \Variables2830[2][0][1] , 
        \Variables2830[4][6][3] , \product1846[4] , \Variables2830[4][2][1] , 
        \Variables2830[4][-4][0] , \TableSelect[3] , \Variables2830[2][4][3] , 
        \Variables2830[2][-7][3] , \Variables2830[0][7][2] , 
        \CycleWaveform34[2] , \Variables2830[1][-7][2] , 
        \Variables2830[1][-3][0] , \TableSelect667[3] , \sum2964[2] , 
        \Variables2830[2][-6][0] , \Variables2830[0][6][1] , Read648, 
        \Variables2830[2][5][0] , OpCodeRegisterWrite, 
        \Variables2830[4][3][2] , \Variables2830[4][-5][3] , 
        \Variables2830[4][7][0] , \Variables2830[4][-1][1] , 
        \Variables2830[2][-2][2] , \Variables2830[2][1][2] , 
        \Variables2830[0][2][3] , n_565, \Variables2830[1][-2][3] , 
        \Variables2830[1][-6][1] , \Variables2830[1][4][0] , 
        \Variables2830[0][-6][2] , \Variables2830[3][7][1] , \Answer639[2] , 
        \Interrupt_Index[0] , \Variables2830[0][-2][0] , 
        \Variables2830[3][3][3] , \Variables2830[1][0][2] , n_399, 
        \RegularWriteRegister_Index848[1] , \Variables2830[3][-2][1] , 
        \Variables2830[3][-6][3] , \MemoryPtr3672[4] , 
        \Variables2830[1][1][1] , \Variables2830[0][-3][3] , 
        \Variables2830[3][2][0] , \Variables2830[4][-8][2] , 
        \Variables2830[0][-7][1] , \Variables2830[3][6][2] , 
        \Variables2830[1][5][3] , \Variables2830[3][-7][0] , 
        \InstructionPtr3995[5] , \Variables2830[3][-3][2] , 
        \ClockCycleCount621[2] , \Answer2629[3] , \n696[3] , n_564, 
        \Variables2830[0][0][1] , \Variables2830[2][3][0] , 
        \Variables2830[4][-3][3] , \Variables2830[4][5][2] , 
        \MemoryPtr3672[0] , \Variables2830[4][-7][1] , 
        \Variables2830[4][1][0] , \Variables2830[0][-8][2] , 
        \Variables2830[2][-4][2] , \Variables2830[2][7][2] , 
        \Variables2830[0][4][3] , \Variables2830[3][-8][3] , 
        \Variables2830[1][-4][3] , \Variables2830[0][5][0] , 
        \Variables2830[2][-5][1] , \Variables2830[2][6][1] , 
        \IPRELOAD_Index[1] , \Variables2830[4][-6][2] , 
        \Variables2830[4][0][3] , \Variables2830[4][-2][0] , 
        \Variables2830[4][4][1] , \Variables2830[2][-1][3] , 
        \Variables2830[2][2][3] , ExceptionJump, \Variables2830[0][1][2] , 
        \InstructionPtr3995[1] , \Variables2830[1][-1][2] , 
        \Variables2830[1][-5][0] , IRQEnable, \Variables2830[1][-1][0] , 
        \ClockCycleCount[2] , \Variables2830[1][-5][2] , \n2831[4][7][3] , 
        \Variables2830[2][-5][3] , \Variables2830[2][6][3] , 
        \Variables2830[0][5][2] , \IPRELOAD_Index[3] , 
        \Variables2830[4][-6][0] , \Variables2830[4][0][1] , 
        \Variables2830[4][-2][2] , \Variables2830[4][4][3] , 
        \Variables2830[0][1][0] , \Variables2830[2][-1][1] , 
        \Variables2830[2][2][1] , \InstructionPtr3995[3] , n_726, n_397, 
        \Variables2830[1][-4][1] , \Variables2830[3][-8][1] , n_691, 
        \Variables2830[2][3][2] , \Variables2830[0][0][3] , 
        \Variables2830[4][-3][1] , \Variables2830[4][5][0] , 
        \MemoryPtr3672[2] , \Variables2830[4][-7][3] , 
        \Variables2830[4][1][2] , \Variables2830[0][4][1] , 
        \Variables2830[2][7][0] , \Variables2830[2][-4][0] , 
        \Variables2830[0][-8][0] , \InstructionPtr3995[7] , 
        \Variables2830[3][-7][2] , \Variables2830[3][-3][0] , \Answer2629[1] , 
        Write657, \Variables2830[0][-3][1] , \Variables2830[3][2][2] , 
        \Variables2830[1][1][3] , \Variables2830[4][-8][0] , \sum1105[1] , 
        \Variables2830[0][-7][3] , \Variables2830[1][5][1] , 
        \Variables2830[3][6][0] , \RegularWriteRegister_Index848[3] , 
        \Variables2830[3][-2][3] , \Variables2830[3][-6][1] , 
        \MemoryPtr3672[6] , \Variables2830[0][-6][0] , 
        \Variables2830[3][7][3] , \Variables2830[1][4][2] , \Answer639[0] , 
        \Interrupt_Index[2] , \Variables2830[0][-2][2] , 
        \Variables2830[1][0][0] , \Variables2830[3][3][1] , n6314, n6315, 
        n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
        n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, 
        n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, 
        n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, 
        n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
        n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
        n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, 
        n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, 
        n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, 
        n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, 
        n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, 
        n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, 
        n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, 
        n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, 
        n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, 
        n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, 
        n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, 
        n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, 
        n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, 
        n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, 
        n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, 
        n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, 
        n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, 
        n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, 
        n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, 
        n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, 
        n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, 
        n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, 
        n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
        n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, 
        n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, 
        n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, 
        n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, 
        n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, 
        n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, 
        n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, 
        n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, 
        n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, 
        n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, 
        n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, 
        n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, 
        n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, 
        n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, 
        n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, 
        n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
        n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, 
        n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
        n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
        n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
        n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
        n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, 
        n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, 
        n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
        n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
        n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
        n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
        n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
        n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
        n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, 
        n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
        n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
        n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, 
        n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
        n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
        n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
        n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, 
        n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
        n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
        n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
        n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
        n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, 
        n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, 
        n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, 
        n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
        n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, 
        n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, 
        n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, 
        n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, 
        n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, 
        n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, 
        n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, 
        n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, 
        n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
        n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, 
        n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
        n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, 
        n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, 
        n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, 
        n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, 
        n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, 
        n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, 
        n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, 
        n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, 
        n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, 
        n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, 
        n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, 
        n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, 
        n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, 
        n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, 
        n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, 
        n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, 
        n7326, n7327, n7328, n7329, net108, net109, net110, net111, net112, 
        n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, 
        n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, 
        \add_417/carry[1] , \add_138/carry[2] , \add_138/carry[1] , 
        \gt_236/AEQB[2] , \*cell*469/U144/Z_0 , \*cell*469/U12/Z_0 , 
        \*cell*469/U11/Z_0 , \*cell*469/U10/Z_0 , \*cell*469/U9/Z_0 , 
        \*cell*469/U7/Z_0 , \*cell*469/U6/Z_0 , n7349;
    tri \Variables[1][7][2]_wire , \Variables[3][4][3]_wire , \MemoryPtr[5] , 
        \Variables[2][-3][0]_wire , \Variables[3][0][1]_wire , 
        \Variables[1][3][0]_wire , \Variables[2][-7][2]_wire , 
        \Variables[4][-4][1]_wire , \InstructionPtr[0] , 
        \Variables[1][-7][3]_wire , \Variables[1][-3][1]_wire , 
        \Variables[4][-5][2]_wire , \Variables[1][2][3]_wire , 
        \Variables[3][1][2]_wire , \Variables[2][-6][1]_wire , 
        \Variables[3][5][0]_wire , \Variables[1][6][1]_wire , 
        \Variables[2][-2][3]_wire , \Variables[4][-1][0]_wire , 
        \Variables[1][-2][2]_wire , \Variables[1][-6][0]_wire , 
        \Variables[4][6][0]_wire , \Variables[0][3][3]_wire , 
        \Variables[2][0][2]_wire , \Variables[0][-5][2]_wire , 
        \Variables[0][-1][0]_wire , \Variables[2][4][0]_wire , 
        \Variables[0][7][1]_wire , \Variables[4][2][2]_wire , 
        \InstructionPtr[4] , \Variables[3][-1][1]_wire , \MemoryPtr[1] , 
        \Variables[3][-5][3]_wire , \Variables[4][3][1]_wire , 
        \Variables[0][6][2]_wire , \Variables[2][5][3]_wire , 
        \Variables[0][-4][1]_wire , \Variables[2][1][1]_wire , 
        \Variables[2][-8][1]_wire , \Variables[0][2][0]_wire , 
        \Variables[4][7][3]_wire , \Variables[3][-4][0]_wire , 
        \Variables[1][-8][0]_wire , \Variables[1][-8][2]_wire , 
        \Variables[3][-4][2]_wire , \Variables[4][3][3]_wire , 
        \Variables[2][5][1]_wire , \Variables[0][6][0]_wire , 
        \Variables[2][1][3]_wire , \Variables[0][2][2]_wire , 
        \Variables[2][-8][3]_wire , \Variables[0][-4][3]_wire , 
        \Variables[4][7][1]_wire , \Variables[3][-1][3]_wire , \MemoryPtr[3] , 
        \Variables[3][-5][1]_wire , \Variables[4][6][2]_wire , 
        \Variables[0][-5][0]_wire , \Variables[2][0][0]_wire , 
        \Variables[0][3][1]_wire , \Variables[0][-1][2]_wire , 
        \Variables[0][7][3]_wire , \Variables[2][4][2]_wire , 
        \Variables[4][2][0]_wire , \InstructionPtr[6] , 
        \Variables[1][-2][0]_wire , Write_wire, \Variables[1][-6][2]_wire , 
        \Variables[4][-5][0]_wire , \Variables[3][1][0]_wire , 
        \Variables[1][2][1]_wire , \Variables[2][-6][3]_wire , 
        \Variables[1][6][3]_wire , \Variables[3][5][2]_wire , 
        \Variables[2][-2][1]_wire , \Variables[4][-1][2]_wire , 
        \Variables[1][-7][1]_wire , \InstructionPtr[2] , 
        \Variables[1][-3][3]_wire , \Variables[1][7][0]_wire , 
        \Variables[3][4][1]_wire , \MemoryPtr[7] , \Variables[2][-3][2]_wire , 
        \Variables[1][3][2]_wire , \Variables[3][0][3]_wire , 
        \Variables[2][-7][0]_wire , \Variables[4][-4][3]_wire , 
        \Variables[3][-7][3]_wire , \Variables[3][-3][1]_wire , 
        \Variables[4][0][2]_wire , \Variables[2][6][0]_wire , 
        \Variables[0][-3][0]_wire , \Variables[0][5][1]_wire , 
        \Variables[0][1][3]_wire , \Variables[0][-7][2]_wire , 
        \Variables[2][2][2]_wire , \Variables[4][-8][1]_wire , 
        \Variables[4][4][0]_wire , \Variables[3][-2][2]_wire , \IRQ[3] , 
        \Variables[3][-6][0]_wire , \Variables[4][5][3]_wire , 
        \Variables[0][-6][1]_wire , \Variables[2][3][1]_wire , 
        \Variables[0][0][0]_wire , \Variables[0][4][2]_wire , 
        \Variables[0][-2][3]_wire , \Variables[2][7][3]_wire , 
        \Variables[4][1][1]_wire , \Variables[1][-1][1]_wire , 
        \Variables[1][-5][3]_wire , \Variables[4][-6][1]_wire , 
        \Variables[2][-5][2]_wire , \Variables[3][2][1]_wire , 
        \Variables[1][1][0]_wire , \Variables[2][-1][0]_wire , 
        \Variables[1][5][2]_wire , \Variables[3][6][3]_wire , 
        \Variables[4][-2][3]_wire , \Variables[1][-4][0]_wire , 
        \Variables[3][-8][0]_wire , \Variables[4][-3][0]_wire , 
        \Variables[3][7][0]_wire , \Variables[1][4][1]_wire , 
        \Variables[2][-4][1]_wire , \Variables[0][-8][1]_wire , 
        \Variables[1][0][3]_wire , \Variables[3][3][2]_wire , 
        \Variables[4][-7][2]_wire , \Variables[4][-3][2]_wire , 
        \Variables[1][4][3]_wire , \Variables[3][7][2]_wire , 
        \Variables[0][-8][3]_wire , \Variables[2][-4][3]_wire , 
        \Variables[3][3][0]_wire , \Variables[1][0][1]_wire , 
        \Variables[4][-7][0]_wire , \Variables[3][-8][2]_wire , 
        \Variables[1][-4][2]_wire , \Variables[4][-6][3]_wire , 
        \Variables[2][-5][0]_wire , \Variables[1][1][2]_wire , 
        \Variables[3][2][3]_wire , \Variables[2][-1][2]_wire , 
        \Variables[3][6][1]_wire , \Variables[1][5][0]_wire , 
        \Variables[4][-2][1]_wire , Read_wire, \Variables[1][-1][3]_wire , 
        \Variables[1][-5][1]_wire , \Variables[4][5][1]_wire , 
        \Variables[0][0][2]_wire , \Variables[0][-6][3]_wire , 
        \Variables[2][3][3]_wire , \Variables[2][7][1]_wire , 
        \Variables[0][-2][1]_wire , \Variables[0][4][0]_wire , 
        \Variables[4][1][3]_wire , \Variables[3][-2][0]_wire , \IRQ[1] , 
        \Variables[3][-6][2]_wire , \Variables[4][0][0]_wire , 
        \Variables[0][5][3]_wire , \Variables[0][-3][2]_wire , 
        \Variables[2][6][2]_wire , \Variables[0][-7][0]_wire , 
        \Variables[2][2][0]_wire , \Variables[0][1][1]_wire , 
        \Variables[4][-8][3]_wire , \Variables[4][4][2]_wire , 
        \Variables[3][-7][1]_wire , \Variables[3][-3][3]_wire , 
        \Variables[2][3][2]_wire , \Variables[0][-6][2]_wire , 
        \Variables[0][0][3]_wire , \Variables[4][5][0]_wire , 
        \Variables[4][1][2]_wire , \Variables[0][4][1]_wire , 
        \Variables[0][-2][0]_wire , \Variables[2][7][0]_wire , 
        \Variables[3][-2][1]_wire , \IRQ[0] , \Variables[3][-6][3]_wire , 
        \Variables[2][6][3]_wire , \Variables[0][-3][3]_wire , 
        \Variables[0][5][2]_wire , \Variables[4][0][1]_wire , 
        \Variables[4][-8][2]_wire , \Variables[4][4][3]_wire , 
        \Variables[0][1][0]_wire , \Variables[0][-7][1]_wire , 
        \Variables[2][2][1]_wire , \Variables[3][-7][0]_wire , 
        \Variables[3][-3][2]_wire , \IRQ[4] , \Variables[3][7][3]_wire , 
        \Variables[1][4][2]_wire , \Variables[4][-3][3]_wire , 
        \Variables[4][-7][1]_wire , \Variables[0][-8][2]_wire , 
        \Variables[2][-4][2]_wire , \Variables[1][0][0]_wire , 
        \Variables[3][3][1]_wire , \Variables[1][-4][3]_wire , 
        \Variables[3][-8][3]_wire , \Variables[2][-5][1]_wire , 
        \Variables[3][2][2]_wire , \Variables[1][1][3]_wire , 
        \Variables[4][-6][2]_wire , \Variables[4][-2][0]_wire , 
        \Variables[2][-1][3]_wire , \Variables[1][5][1]_wire , 
        \Variables[3][6][0]_wire , \Variables[1][-1][2]_wire , 
        \Variables[1][-5][0]_wire , \Variables[1][-1][0]_wire , 
        \Variables[1][-5][2]_wire , \Variables[2][-5][3]_wire , 
        \Variables[1][1][1]_wire , \Variables[3][2][0]_wire , 
        \Variables[4][-6][0]_wire , \Variables[4][-2][2]_wire , 
        \Variables[2][-1][1]_wire , \Variables[3][6][2]_wire , 
        \Variables[1][5][3]_wire , \Variables[1][-4][1]_wire , 
        \Variables[3][-8][1]_wire , \Variables[1][4][0]_wire , 
        \Variables[3][7][1]_wire , \Variables[4][-3][1]_wire , 
        \Variables[4][-7][3]_wire , \Variables[2][-4][0]_wire , 
        \Variables[0][-8][0]_wire , \Variables[3][3][3]_wire , 
        \Variables[1][0][2]_wire , \Variables[3][-7][2]_wire , 
        \Variables[3][-3][0]_wire , \Variables[0][5][0]_wire , 
        \Variables[0][-3][1]_wire , \Variables[2][6][1]_wire , 
        \Variables[4][0][3]_wire , \Variables[4][-8][0]_wire , 
        \Variables[4][4][1]_wire , \Variables[0][-7][3]_wire , 
        \Variables[2][2][3]_wire , \Variables[0][1][2]_wire , 
        \Variables[3][-2][3]_wire , \Variables[3][-6][1]_wire , \IRQ[2] , 
        \Variables[0][0][1]_wire , \Variables[0][-6][0]_wire , 
        \Variables[2][3][0]_wire , \Variables[4][5][2]_wire , 
        \Variables[4][1][0]_wire , \Variables[2][7][2]_wire , 
        \Variables[0][-2][2]_wire , \Variables[0][4][3]_wire , 
        \Variables[1][-2][1]_wire , \Variables[1][-6][3]_wire , 
        \Variables[1][2][0]_wire , \Variables[3][1][1]_wire , 
        \Variables[2][-6][2]_wire , \Variables[4][-5][1]_wire , 
        \Variables[4][-1][3]_wire , \Variables[3][5][3]_wire , 
        \Variables[1][6][2]_wire , \Variables[2][-2][0]_wire , 
        \InstructionPtr[3] , \Variables[1][-7][0]_wire , 
        \Variables[1][-3][2]_wire , \Variables[1][7][1]_wire , 
        \Variables[3][4][0]_wire , \MemoryPtr[6] , \Variables[2][-3][3]_wire , 
        \Variables[4][-4][2]_wire , \Variables[3][0][2]_wire , 
        \Variables[1][3][3]_wire , \Variables[2][-7][1]_wire , 
        \Variables[1][-8][3]_wire , \Variables[3][-4][3]_wire , 
        \Variables[0][6][1]_wire , \Variables[2][5][0]_wire , 
        \Variables[4][3][2]_wire , \Variables[4][7][0]_wire , 
        \Variables[0][-4][2]_wire , \Variables[2][-8][2]_wire , 
        \Variables[2][1][2]_wire , \Variables[0][2][3]_wire , 
        \Variables[3][-1][2]_wire , \Variables[3][-5][0]_wire , \MemoryPtr[2] , 
        \Variables[0][3][0]_wire , \Variables[2][0][1]_wire , 
        \Variables[0][-5][1]_wire , \Variables[4][2][1]_wire , 
        \Variables[4][6][3]_wire , \InstructionPtr[7] , 
        \Variables[0][-1][3]_wire , \Variables[0][7][2]_wire , 
        \Variables[2][4][3]_wire , \Variables[0][-5][3]_wire , 
        \Variables[2][0][3]_wire , \Variables[0][3][2]_wire , 
        \Variables[4][6][1]_wire , \Variables[4][2][3]_wire , 
        \InstructionPtr[5] , \Variables[0][-1][1]_wire , 
        \Variables[0][7][0]_wire , \Variables[2][4][1]_wire , 
        \Variables[3][-1][0]_wire , \Variables[3][-5][2]_wire , \MemoryPtr[0] , 
        \Variables[2][5][2]_wire , \Variables[0][6][3]_wire , 
        \Variables[4][3][0]_wire , \Variables[4][7][2]_wire , 
        \Variables[0][2][1]_wire , \Variables[2][1][0]_wire , 
        \Variables[0][-4][0]_wire , \Variables[2][-8][0]_wire , 
        \Variables[3][-4][1]_wire , \Variables[1][-8][1]_wire , 
        \Variables[3][4][2]_wire , \MemoryPtr[4] , \Variables[1][7][3]_wire , 
        \Variables[2][-3][1]_wire , \Variables[4][-4][0]_wire , 
        \Variables[1][3][1]_wire , \Variables[3][0][0]_wire , 
        \Variables[2][-7][3]_wire , \Variables[1][-7][2]_wire , 
        \InstructionPtr[1] , \Variables[1][-3][0]_wire , 
        \Variables[3][1][3]_wire , \Variables[1][2][2]_wire , 
        \Variables[2][-6][0]_wire , \Variables[4][-5][3]_wire , 
        \Variables[4][-1][1]_wire , \Variables[1][6][0]_wire , 
        \Variables[3][5][1]_wire , \Variables[2][-2][2]_wire , 
        \Variables[1][-2][3]_wire , \Variables[1][-6][1]_wire ;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 , SYNOPSYS_UNCONNECTED_4 ;
    tran( \Variables[0][-8][3]_wire , \Variables[0][-8][3]  );
    tran( \Variables[0][-8][2]_wire , \Variables[0][-8][2]  );
    tran( \Variables[0][-8][1]_wire , \Variables[0][-8][1]  );
    tran( \Variables[0][-8][0]_wire , \Variables[0][-8][0]  );
    tran( \Variables[0][-7][3]_wire , \Variables[0][-7][3]  );
    tran( \Variables[0][-7][2]_wire , \Variables[0][-7][2]  );
    tran( \Variables[0][-7][1]_wire , \Variables[0][-7][1]  );
    tran( \Variables[0][-7][0]_wire , \Variables[0][-7][0]  );
    tran( \Variables[0][-6][3]_wire , \Variables[0][-6][3]  );
    tran( \Variables[0][-6][2]_wire , \Variables[0][-6][2]  );
    tran( \Variables[0][-6][1]_wire , \Variables[0][-6][1]  );
    tran( \Variables[0][-6][0]_wire , \Variables[0][-6][0]  );
    tran( \Variables[0][-5][3]_wire , \Variables[0][-5][3]  );
    tran( \Variables[0][-5][2]_wire , \Variables[0][-5][2]  );
    tran( \Variables[0][-5][1]_wire , \Variables[0][-5][1]  );
    tran( \Variables[0][-5][0]_wire , \Variables[0][-5][0]  );
    tran( \Variables[0][-4][3]_wire , \Variables[0][-4][3]  );
    tran( \Variables[0][-4][2]_wire , \Variables[0][-4][2]  );
    tran( \Variables[0][-4][1]_wire , \Variables[0][-4][1]  );
    tran( \Variables[0][-4][0]_wire , \Variables[0][-4][0]  );
    tran( \Variables[0][-3][3]_wire , \Variables[0][-3][3]  );
    tran( \Variables[0][-3][2]_wire , \Variables[0][-3][2]  );
    tran( \Variables[0][-3][1]_wire , \Variables[0][-3][1]  );
    tran( \Variables[0][-3][0]_wire , \Variables[0][-3][0]  );
    tran( \Variables[0][-2][3]_wire , \Variables[0][-2][3]  );
    tran( \Variables[0][-2][2]_wire , \Variables[0][-2][2]  );
    tran( \Variables[0][-2][1]_wire , \Variables[0][-2][1]  );
    tran( \Variables[0][-2][0]_wire , \Variables[0][-2][0]  );
    tran( \Variables[0][-1][3]_wire , \Variables[0][-1][3]  );
    tran( \Variables[0][-1][2]_wire , \Variables[0][-1][2]  );
    tran( \Variables[0][-1][1]_wire , \Variables[0][-1][1]  );
    tran( \Variables[0][-1][0]_wire , \Variables[0][-1][0]  );
    tran( \Variables[0][0][3]_wire , \Variables[0][0][3]  );
    tran( \Variables[0][0][2]_wire , \Variables[0][0][2]  );
    tran( \Variables[0][0][1]_wire , \Variables[0][0][1]  );
    tran( \Variables[0][0][0]_wire , \Variables[0][0][0]  );
    tran( \Variables[0][1][3]_wire , \Variables[0][1][3]  );
    tran( \Variables[0][1][2]_wire , \Variables[0][1][2]  );
    tran( \Variables[0][1][1]_wire , \Variables[0][1][1]  );
    tran( \Variables[0][1][0]_wire , \Variables[0][1][0]  );
    tran( \Variables[0][2][3]_wire , \Variables[0][2][3]  );
    tran( \Variables[0][2][2]_wire , \Variables[0][2][2]  );
    tran( \Variables[0][2][1]_wire , \Variables[0][2][1]  );
    tran( \Variables[0][2][0]_wire , \Variables[0][2][0]  );
    tran( \Variables[0][3][3]_wire , \Variables[0][3][3]  );
    tran( \Variables[0][3][2]_wire , \Variables[0][3][2]  );
    tran( \Variables[0][3][1]_wire , \Variables[0][3][1]  );
    tran( \Variables[0][3][0]_wire , \Variables[0][3][0]  );
    tran( \Variables[0][4][3]_wire , \Variables[0][4][3]  );
    tran( \Variables[0][4][2]_wire , \Variables[0][4][2]  );
    tran( \Variables[0][4][1]_wire , \Variables[0][4][1]  );
    tran( \Variables[0][4][0]_wire , \Variables[0][4][0]  );
    tran( \Variables[0][5][3]_wire , \Variables[0][5][3]  );
    tran( \Variables[0][5][2]_wire , \Variables[0][5][2]  );
    tran( \Variables[0][5][1]_wire , \Variables[0][5][1]  );
    tran( \Variables[0][5][0]_wire , \Variables[0][5][0]  );
    tran( \Variables[0][6][3]_wire , \Variables[0][6][3]  );
    tran( \Variables[0][6][2]_wire , \Variables[0][6][2]  );
    tran( \Variables[0][6][1]_wire , \Variables[0][6][1]  );
    tran( \Variables[0][6][0]_wire , \Variables[0][6][0]  );
    tran( \Variables[0][7][3]_wire , \Variables[0][7][3]  );
    tran( \Variables[0][7][2]_wire , \Variables[0][7][2]  );
    tran( \Variables[0][7][1]_wire , \Variables[0][7][1]  );
    tran( \Variables[0][7][0]_wire , \Variables[0][7][0]  );
    tran( \Variables[1][-8][3]_wire , \Variables[1][-8][3]  );
    tran( \Variables[1][-8][2]_wire , \Variables[1][-8][2]  );
    tran( \Variables[1][-8][1]_wire , \Variables[1][-8][1]  );
    tran( \Variables[1][-8][0]_wire , \Variables[1][-8][0]  );
    tran( \Variables[1][-7][3]_wire , \Variables[1][-7][3]  );
    tran( \Variables[1][-7][2]_wire , \Variables[1][-7][2]  );
    tran( \Variables[1][-7][1]_wire , \Variables[1][-7][1]  );
    tran( \Variables[1][-7][0]_wire , \Variables[1][-7][0]  );
    tran( \Variables[1][-6][3]_wire , \Variables[1][-6][3]  );
    tran( \Variables[1][-6][2]_wire , \Variables[1][-6][2]  );
    tran( \Variables[1][-6][1]_wire , \Variables[1][-6][1]  );
    tran( \Variables[1][-6][0]_wire , \Variables[1][-6][0]  );
    tran( \Variables[1][-5][3]_wire , \Variables[1][-5][3]  );
    tran( \Variables[1][-5][2]_wire , \Variables[1][-5][2]  );
    tran( \Variables[1][-5][1]_wire , \Variables[1][-5][1]  );
    tran( \Variables[1][-5][0]_wire , \Variables[1][-5][0]  );
    tran( \Variables[1][-4][3]_wire , \Variables[1][-4][3]  );
    tran( \Variables[1][-4][2]_wire , \Variables[1][-4][2]  );
    tran( \Variables[1][-4][1]_wire , \Variables[1][-4][1]  );
    tran( \Variables[1][-4][0]_wire , \Variables[1][-4][0]  );
    tran( \Variables[1][-3][3]_wire , \Variables[1][-3][3]  );
    tran( \Variables[1][-3][2]_wire , \Variables[1][-3][2]  );
    tran( \Variables[1][-3][1]_wire , \Variables[1][-3][1]  );
    tran( \Variables[1][-3][0]_wire , \Variables[1][-3][0]  );
    tran( \Variables[1][-2][3]_wire , \Variables[1][-2][3]  );
    tran( \Variables[1][-2][2]_wire , \Variables[1][-2][2]  );
    tran( \Variables[1][-2][1]_wire , \Variables[1][-2][1]  );
    tran( \Variables[1][-2][0]_wire , \Variables[1][-2][0]  );
    tran( \Variables[1][-1][3]_wire , \Variables[1][-1][3]  );
    tran( \Variables[1][-1][2]_wire , \Variables[1][-1][2]  );
    tran( \Variables[1][-1][1]_wire , \Variables[1][-1][1]  );
    tran( \Variables[1][-1][0]_wire , \Variables[1][-1][0]  );
    tran( \Variables[1][0][3]_wire , \Variables[1][0][3]  );
    tran( \Variables[1][0][2]_wire , \Variables[1][0][2]  );
    tran( \Variables[1][0][1]_wire , \Variables[1][0][1]  );
    tran( \Variables[1][0][0]_wire , \Variables[1][0][0]  );
    tran( \Variables[1][1][3]_wire , \Variables[1][1][3]  );
    tran( \Variables[1][1][2]_wire , \Variables[1][1][2]  );
    tran( \Variables[1][1][1]_wire , \Variables[1][1][1]  );
    tran( \Variables[1][1][0]_wire , \Variables[1][1][0]  );
    tran( \Variables[1][2][3]_wire , \Variables[1][2][3]  );
    tran( \Variables[1][2][2]_wire , \Variables[1][2][2]  );
    tran( \Variables[1][2][1]_wire , \Variables[1][2][1]  );
    tran( \Variables[1][2][0]_wire , \Variables[1][2][0]  );
    tran( \Variables[1][3][3]_wire , \Variables[1][3][3]  );
    tran( \Variables[1][3][2]_wire , \Variables[1][3][2]  );
    tran( \Variables[1][3][1]_wire , \Variables[1][3][1]  );
    tran( \Variables[1][3][0]_wire , \Variables[1][3][0]  );
    tran( \Variables[1][4][3]_wire , \Variables[1][4][3]  );
    tran( \Variables[1][4][2]_wire , \Variables[1][4][2]  );
    tran( \Variables[1][4][1]_wire , \Variables[1][4][1]  );
    tran( \Variables[1][4][0]_wire , \Variables[1][4][0]  );
    tran( \Variables[1][5][3]_wire , \Variables[1][5][3]  );
    tran( \Variables[1][5][2]_wire , \Variables[1][5][2]  );
    tran( \Variables[1][5][1]_wire , \Variables[1][5][1]  );
    tran( \Variables[1][5][0]_wire , \Variables[1][5][0]  );
    tran( \Variables[1][6][3]_wire , \Variables[1][6][3]  );
    tran( \Variables[1][6][2]_wire , \Variables[1][6][2]  );
    tran( \Variables[1][6][1]_wire , \Variables[1][6][1]  );
    tran( \Variables[1][6][0]_wire , \Variables[1][6][0]  );
    tran( \Variables[1][7][3]_wire , \Variables[1][7][3]  );
    tran( \Variables[1][7][2]_wire , \Variables[1][7][2]  );
    tran( \Variables[1][7][1]_wire , \Variables[1][7][1]  );
    tran( \Variables[1][7][0]_wire , \Variables[1][7][0]  );
    tran( \Variables[2][-8][3]_wire , \Variables[2][-8][3]  );
    tran( \Variables[2][-8][2]_wire , \Variables[2][-8][2]  );
    tran( \Variables[2][-8][1]_wire , \Variables[2][-8][1]  );
    tran( \Variables[2][-8][0]_wire , \Variables[2][-8][0]  );
    tran( \Variables[2][-7][3]_wire , \Variables[2][-7][3]  );
    tran( \Variables[2][-7][2]_wire , \Variables[2][-7][2]  );
    tran( \Variables[2][-7][1]_wire , \Variables[2][-7][1]  );
    tran( \Variables[2][-7][0]_wire , \Variables[2][-7][0]  );
    tran( \Variables[2][-6][3]_wire , \Variables[2][-6][3]  );
    tran( \Variables[2][-6][2]_wire , \Variables[2][-6][2]  );
    tran( \Variables[2][-6][1]_wire , \Variables[2][-6][1]  );
    tran( \Variables[2][-6][0]_wire , \Variables[2][-6][0]  );
    tran( \Variables[2][-5][3]_wire , \Variables[2][-5][3]  );
    tran( \Variables[2][-5][2]_wire , \Variables[2][-5][2]  );
    tran( \Variables[2][-5][1]_wire , \Variables[2][-5][1]  );
    tran( \Variables[2][-5][0]_wire , \Variables[2][-5][0]  );
    tran( \Variables[2][-4][3]_wire , \Variables[2][-4][3]  );
    tran( \Variables[2][-4][2]_wire , \Variables[2][-4][2]  );
    tran( \Variables[2][-4][1]_wire , \Variables[2][-4][1]  );
    tran( \Variables[2][-4][0]_wire , \Variables[2][-4][0]  );
    tran( \Variables[2][-3][3]_wire , \Variables[2][-3][3]  );
    tran( \Variables[2][-3][2]_wire , \Variables[2][-3][2]  );
    tran( \Variables[2][-3][1]_wire , \Variables[2][-3][1]  );
    tran( \Variables[2][-3][0]_wire , \Variables[2][-3][0]  );
    tran( \Variables[2][-2][3]_wire , \Variables[2][-2][3]  );
    tran( \Variables[2][-2][2]_wire , \Variables[2][-2][2]  );
    tran( \Variables[2][-2][1]_wire , \Variables[2][-2][1]  );
    tran( \Variables[2][-2][0]_wire , \Variables[2][-2][0]  );
    tran( \Variables[2][-1][3]_wire , \Variables[2][-1][3]  );
    tran( \Variables[2][-1][2]_wire , \Variables[2][-1][2]  );
    tran( \Variables[2][-1][1]_wire , \Variables[2][-1][1]  );
    tran( \Variables[2][-1][0]_wire , \Variables[2][-1][0]  );
    tran( \Variables[2][0][3]_wire , \Variables[2][0][3]  );
    tran( \Variables[2][0][2]_wire , \Variables[2][0][2]  );
    tran( \Variables[2][0][1]_wire , \Variables[2][0][1]  );
    tran( \Variables[2][0][0]_wire , \Variables[2][0][0]  );
    tran( \Variables[2][1][3]_wire , \Variables[2][1][3]  );
    tran( \Variables[2][1][2]_wire , \Variables[2][1][2]  );
    tran( \Variables[2][1][1]_wire , \Variables[2][1][1]  );
    tran( \Variables[2][1][0]_wire , \Variables[2][1][0]  );
    tran( \Variables[2][2][3]_wire , \Variables[2][2][3]  );
    tran( \Variables[2][2][2]_wire , \Variables[2][2][2]  );
    tran( \Variables[2][2][1]_wire , \Variables[2][2][1]  );
    tran( \Variables[2][2][0]_wire , \Variables[2][2][0]  );
    tran( \Variables[2][3][3]_wire , \Variables[2][3][3]  );
    tran( \Variables[2][3][2]_wire , \Variables[2][3][2]  );
    tran( \Variables[2][3][1]_wire , \Variables[2][3][1]  );
    tran( \Variables[2][3][0]_wire , \Variables[2][3][0]  );
    tran( \Variables[2][4][3]_wire , \Variables[2][4][3]  );
    tran( \Variables[2][4][2]_wire , \Variables[2][4][2]  );
    tran( \Variables[2][4][1]_wire , \Variables[2][4][1]  );
    tran( \Variables[2][4][0]_wire , \Variables[2][4][0]  );
    tran( \Variables[2][5][3]_wire , \Variables[2][5][3]  );
    tran( \Variables[2][5][2]_wire , \Variables[2][5][2]  );
    tran( \Variables[2][5][1]_wire , \Variables[2][5][1]  );
    tran( \Variables[2][5][0]_wire , \Variables[2][5][0]  );
    tran( \Variables[2][6][3]_wire , \Variables[2][6][3]  );
    tran( \Variables[2][6][2]_wire , \Variables[2][6][2]  );
    tran( \Variables[2][6][1]_wire , \Variables[2][6][1]  );
    tran( \Variables[2][6][0]_wire , \Variables[2][6][0]  );
    tran( \Variables[2][7][3]_wire , \Variables[2][7][3]  );
    tran( \Variables[2][7][2]_wire , \Variables[2][7][2]  );
    tran( \Variables[2][7][1]_wire , \Variables[2][7][1]  );
    tran( \Variables[2][7][0]_wire , \Variables[2][7][0]  );
    tran( \Variables[3][-8][3]_wire , \Variables[3][-8][3]  );
    tran( \Variables[3][-8][2]_wire , \Variables[3][-8][2]  );
    tran( \Variables[3][-8][1]_wire , \Variables[3][-8][1]  );
    tran( \Variables[3][-8][0]_wire , \Variables[3][-8][0]  );
    tran( \Variables[3][-7][3]_wire , \Variables[3][-7][3]  );
    tran( \Variables[3][-7][2]_wire , \Variables[3][-7][2]  );
    tran( \Variables[3][-7][1]_wire , \Variables[3][-7][1]  );
    tran( \Variables[3][-7][0]_wire , \Variables[3][-7][0]  );
    tran( \Variables[3][-6][3]_wire , \Variables[3][-6][3]  );
    tran( \Variables[3][-6][2]_wire , \Variables[3][-6][2]  );
    tran( \Variables[3][-6][1]_wire , \Variables[3][-6][1]  );
    tran( \Variables[3][-6][0]_wire , \Variables[3][-6][0]  );
    tran( \Variables[3][-5][3]_wire , \Variables[3][-5][3]  );
    tran( \Variables[3][-5][2]_wire , \Variables[3][-5][2]  );
    tran( \Variables[3][-5][1]_wire , \Variables[3][-5][1]  );
    tran( \Variables[3][-5][0]_wire , \Variables[3][-5][0]  );
    tran( \Variables[3][-4][3]_wire , \Variables[3][-4][3]  );
    tran( \Variables[3][-4][2]_wire , \Variables[3][-4][2]  );
    tran( \Variables[3][-4][1]_wire , \Variables[3][-4][1]  );
    tran( \Variables[3][-4][0]_wire , \Variables[3][-4][0]  );
    tran( \Variables[3][-3][3]_wire , \Variables[3][-3][3]  );
    tran( \Variables[3][-3][2]_wire , \Variables[3][-3][2]  );
    tran( \Variables[3][-3][1]_wire , \Variables[3][-3][1]  );
    tran( \Variables[3][-3][0]_wire , \Variables[3][-3][0]  );
    tran( \Variables[3][-2][3]_wire , \Variables[3][-2][3]  );
    tran( \Variables[3][-2][2]_wire , \Variables[3][-2][2]  );
    tran( \Variables[3][-2][1]_wire , \Variables[3][-2][1]  );
    tran( \Variables[3][-2][0]_wire , \Variables[3][-2][0]  );
    tran( \Variables[3][-1][3]_wire , \Variables[3][-1][3]  );
    tran( \Variables[3][-1][2]_wire , \Variables[3][-1][2]  );
    tran( \Variables[3][-1][1]_wire , \Variables[3][-1][1]  );
    tran( \Variables[3][-1][0]_wire , \Variables[3][-1][0]  );
    tran( \Variables[3][0][3]_wire , \Variables[3][0][3]  );
    tran( \Variables[3][0][2]_wire , \Variables[3][0][2]  );
    tran( \Variables[3][0][1]_wire , \Variables[3][0][1]  );
    tran( \Variables[3][0][0]_wire , \Variables[3][0][0]  );
    tran( \Variables[3][1][3]_wire , \Variables[3][1][3]  );
    tran( \Variables[3][1][2]_wire , \Variables[3][1][2]  );
    tran( \Variables[3][1][1]_wire , \Variables[3][1][1]  );
    tran( \Variables[3][1][0]_wire , \Variables[3][1][0]  );
    tran( \Variables[3][2][3]_wire , \Variables[3][2][3]  );
    tran( \Variables[3][2][2]_wire , \Variables[3][2][2]  );
    tran( \Variables[3][2][1]_wire , \Variables[3][2][1]  );
    tran( \Variables[3][2][0]_wire , \Variables[3][2][0]  );
    tran( \Variables[3][3][3]_wire , \Variables[3][3][3]  );
    tran( \Variables[3][3][2]_wire , \Variables[3][3][2]  );
    tran( \Variables[3][3][1]_wire , \Variables[3][3][1]  );
    tran( \Variables[3][3][0]_wire , \Variables[3][3][0]  );
    tran( \Variables[3][4][3]_wire , \Variables[3][4][3]  );
    tran( \Variables[3][4][2]_wire , \Variables[3][4][2]  );
    tran( \Variables[3][4][1]_wire , \Variables[3][4][1]  );
    tran( \Variables[3][4][0]_wire , \Variables[3][4][0]  );
    tran( \Variables[3][5][3]_wire , \Variables[3][5][3]  );
    tran( \Variables[3][5][2]_wire , \Variables[3][5][2]  );
    tran( \Variables[3][5][1]_wire , \Variables[3][5][1]  );
    tran( \Variables[3][5][0]_wire , \Variables[3][5][0]  );
    tran( \Variables[3][6][3]_wire , \Variables[3][6][3]  );
    tran( \Variables[3][6][2]_wire , \Variables[3][6][2]  );
    tran( \Variables[3][6][1]_wire , \Variables[3][6][1]  );
    tran( \Variables[3][6][0]_wire , \Variables[3][6][0]  );
    tran( \Variables[3][7][3]_wire , \Variables[3][7][3]  );
    tran( \Variables[3][7][2]_wire , \Variables[3][7][2]  );
    tran( \Variables[3][7][1]_wire , \Variables[3][7][1]  );
    tran( \Variables[3][7][0]_wire , \Variables[3][7][0]  );
    tran( \Variables[4][-8][3]_wire , \Variables[4][-8][3]  );
    tran( \Variables[4][-8][2]_wire , \Variables[4][-8][2]  );
    tran( \Variables[4][-8][1]_wire , \Variables[4][-8][1]  );
    tran( \Variables[4][-8][0]_wire , \Variables[4][-8][0]  );
    tran( \Variables[4][-7][3]_wire , \Variables[4][-7][3]  );
    tran( \Variables[4][-7][2]_wire , \Variables[4][-7][2]  );
    tran( \Variables[4][-7][1]_wire , \Variables[4][-7][1]  );
    tran( \Variables[4][-7][0]_wire , \Variables[4][-7][0]  );
    tran( \Variables[4][-6][3]_wire , \Variables[4][-6][3]  );
    tran( \Variables[4][-6][2]_wire , \Variables[4][-6][2]  );
    tran( \Variables[4][-6][1]_wire , \Variables[4][-6][1]  );
    tran( \Variables[4][-6][0]_wire , \Variables[4][-6][0]  );
    tran( \Variables[4][-5][3]_wire , \Variables[4][-5][3]  );
    tran( \Variables[4][-5][2]_wire , \Variables[4][-5][2]  );
    tran( \Variables[4][-5][1]_wire , \Variables[4][-5][1]  );
    tran( \Variables[4][-5][0]_wire , \Variables[4][-5][0]  );
    tran( \Variables[4][-4][3]_wire , \Variables[4][-4][3]  );
    tran( \Variables[4][-4][2]_wire , \Variables[4][-4][2]  );
    tran( \Variables[4][-4][1]_wire , \Variables[4][-4][1]  );
    tran( \Variables[4][-4][0]_wire , \Variables[4][-4][0]  );
    tran( \Variables[4][-3][3]_wire , \Variables[4][-3][3]  );
    tran( \Variables[4][-3][2]_wire , \Variables[4][-3][2]  );
    tran( \Variables[4][-3][1]_wire , \Variables[4][-3][1]  );
    tran( \Variables[4][-3][0]_wire , \Variables[4][-3][0]  );
    tran( \Variables[4][-2][3]_wire , \Variables[4][-2][3]  );
    tran( \Variables[4][-2][2]_wire , \Variables[4][-2][2]  );
    tran( \Variables[4][-2][1]_wire , \Variables[4][-2][1]  );
    tran( \Variables[4][-2][0]_wire , \Variables[4][-2][0]  );
    tran( \Variables[4][-1][3]_wire , \Variables[4][-1][3]  );
    tran( \Variables[4][-1][2]_wire , \Variables[4][-1][2]  );
    tran( \Variables[4][-1][1]_wire , \Variables[4][-1][1]  );
    tran( \Variables[4][-1][0]_wire , \Variables[4][-1][0]  );
    tran( \Variables[4][0][3]_wire , \Variables[4][0][3]  );
    tran( \Variables[4][0][2]_wire , \Variables[4][0][2]  );
    tran( \Variables[4][0][1]_wire , \Variables[4][0][1]  );
    tran( \Variables[4][0][0]_wire , \Variables[4][0][0]  );
    tran( \Variables[4][1][3]_wire , \Variables[4][1][3]  );
    tran( \Variables[4][1][2]_wire , \Variables[4][1][2]  );
    tran( \Variables[4][1][1]_wire , \Variables[4][1][1]  );
    tran( \Variables[4][1][0]_wire , \Variables[4][1][0]  );
    tran( \Variables[4][2][3]_wire , \Variables[4][2][3]  );
    tran( \Variables[4][2][2]_wire , \Variables[4][2][2]  );
    tran( \Variables[4][2][1]_wire , \Variables[4][2][1]  );
    tran( \Variables[4][2][0]_wire , \Variables[4][2][0]  );
    tran( \Variables[4][3][3]_wire , \Variables[4][3][3]  );
    tran( \Variables[4][3][2]_wire , \Variables[4][3][2]  );
    tran( \Variables[4][3][1]_wire , \Variables[4][3][1]  );
    tran( \Variables[4][3][0]_wire , \Variables[4][3][0]  );
    tran( \Variables[4][4][3]_wire , \Variables[4][4][3]  );
    tran( \Variables[4][4][2]_wire , \Variables[4][4][2]  );
    tran( \Variables[4][4][1]_wire , \Variables[4][4][1]  );
    tran( \Variables[4][4][0]_wire , \Variables[4][4][0]  );
    tran( \Variables[4][5][3]_wire , \Variables[4][5][3]  );
    tran( \Variables[4][5][2]_wire , \Variables[4][5][2]  );
    tran( \Variables[4][5][1]_wire , \Variables[4][5][1]  );
    tran( \Variables[4][5][0]_wire , \Variables[4][5][0]  );
    tran( \Variables[4][6][3]_wire , \Variables[4][6][3]  );
    tran( \Variables[4][6][2]_wire , \Variables[4][6][2]  );
    tran( \Variables[4][6][1]_wire , \Variables[4][6][1]  );
    tran( \Variables[4][6][0]_wire , \Variables[4][6][0]  );
    tran( \Variables[4][7][3]_wire , \Variables[4][7][3]  );
    tran( \Variables[4][7][2]_wire , \Variables[4][7][2]  );
    tran( \Variables[4][7][1]_wire , \Variables[4][7][1]  );
    tran( \Variables[4][7][0]_wire , \Variables[4][7][0]  );
    tran( \InstructionPtr[7] , InstructionPtr[7] );
    tran( \InstructionPtr[6] , InstructionPtr[6] );
    tran( \InstructionPtr[5] , InstructionPtr[5] );
    tran( \InstructionPtr[4] , InstructionPtr[4] );
    tran( \InstructionPtr[3] , InstructionPtr[3] );
    tran( \InstructionPtr[2] , InstructionPtr[2] );
    tran( \InstructionPtr[1] , InstructionPtr[1] );
    tran( \InstructionPtr[0] , InstructionPtr[0] );
    tran( \MemoryPtr[7] , MemoryPtr[7] );
    tran( \MemoryPtr[6] , MemoryPtr[6] );
    tran( \MemoryPtr[5] , MemoryPtr[5] );
    tran( \MemoryPtr[4] , MemoryPtr[4] );
    tran( \MemoryPtr[3] , MemoryPtr[3] );
    tran( \MemoryPtr[2] , MemoryPtr[2] );
    tran( \MemoryPtr[1] , MemoryPtr[1] );
    tran( \MemoryPtr[0] , MemoryPtr[0] );
    tran( Read_wire, Read );
    tran( Write_wire, Write );
    tran( \IRQ[0] , IRQ[0] );
    tran( \IRQ[1] , IRQ[1] );
    tran( \IRQ[2] , IRQ[2] );
    tran( \IRQ[3] , IRQ[3] );
    tran( \IRQ[4] , IRQ[4] );
    GTECH_ZERO U1110 ( .Z(n7348) );
    GTECH_ONE U1111 ( .Z(n7349) );
    GTECH_OAI2N2 U1112 ( .A(n6314), .B(\add_138/carry[2] ), .C(n6314), .D(
        \add_138/carry[2] ), .Z(\sum1105[2] ) );
    GTECH_NOT U1113 ( .A(\ClockCycleCount[2] ), .Z(n6314) );
    GTECH_AND_NOT U1114 ( .A(\ClockCycleCount[1] ), .B(n6315), .Z(
        \add_138/carry[2] ) );
    GTECH_OAI2N2 U1115 ( .A(\ClockCycleCount[1] ), .B(n6315), .C(
        \ClockCycleCount[1] ), .D(n6315), .Z(\sum1105[1] ) );
    GTECH_NOT U1116 ( .A(\add_138/carry[1] ), .Z(n6315) );
    GTECH_NOT U1117 ( .A(\add_138/carry[1] ), .Z(\sum1105[0] ) );
    GTECH_OR_NOT U1118 ( .A(\TableSelect[3] ), .B(n6316), .Z(
        OutOfRangeException2645) );
    GTECH_OR_NOT U1119 ( .A(Read_wire), .B(n6317), .Z(\n3651[7] ) );
    GTECH_OR2 U1120 ( .A(ExceptionJump), .B(n6318), .Z(n_4166) );
    GTECH_NAND2 U1121 ( .A(n6319), .B(\IRQ2736[4] ), .Z(n_693) );
    GTECH_OAI21 U1122 ( .A(n6320), .B(n6321), .C(n6322), .Z(n_692) );
    GTECH_OAI21 U1123 ( .A(n6320), .B(n6323), .C(n6322), .Z(n_691) );
    GTECH_NAND2 U1124 ( .A(n6322), .B(n6324), .Z(n_690) );
    GTECH_OAI21 U1125 ( .A(n6320), .B(n6325), .C(n6322), .Z(n_689) );
    GTECH_AND2 U1126 ( .A(n6322), .B(n_660), .Z(n_726) );
    GTECH_OA21 U1127 ( .A(n6326), .B(n6327), .C(n6328), .Z(\*cell*469/U6/Z_0 )
         );
    GTECH_AO21 U1128 ( .A(n6329), .B(n6330), .C(\*cell*469/U12/Z_0 ), .Z(
        \*cell*469/U9/Z_0 ) );
    GTECH_AO22 U1129 ( .A(n6328), .B(n6331), .C(n6329), .D(n6332), .Z(
        \*cell*469/U10/Z_0 ) );
    GTECH_AND2 U1130 ( .A(n6333), .B(n6334), .Z(\*cell*469/U11/Z_0 ) );
    GTECH_AND2 U1131 ( .A(n6336), .B(\Upper[3] ), .Z(n6335) );
    GTECH_NOT U1132 ( .A(n6337), .Z(\Variables2830[0][-8][3] ) );
    GTECH_NOT U1133 ( .A(n6338), .Z(\Variables2830[0][-8][2] ) );
    GTECH_NOT U1134 ( .A(n6339), .Z(\Variables2830[0][-8][1] ) );
    GTECH_NOT U1135 ( .A(n6340), .Z(\Variables2830[0][-8][0] ) );
    GTECH_NOT U1136 ( .A(n6341), .Z(\Variables2830[0][-7][3] ) );
    GTECH_NOT U1137 ( .A(n6342), .Z(\Variables2830[0][-7][2] ) );
    GTECH_NOT U1138 ( .A(n6343), .Z(\Variables2830[0][-7][1] ) );
    GTECH_NOT U1139 ( .A(n6344), .Z(\Variables2830[0][-7][0] ) );
    GTECH_OAI2N2 U1140 ( .A(n6345), .B(n6346), .C(\Variables[0][-6][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-6][3] ) );
    GTECH_OAI2N2 U1141 ( .A(n6348), .B(n6346), .C(\Variables[0][-6][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-6][2] ) );
    GTECH_OAI2N2 U1142 ( .A(n6349), .B(n6346), .C(\Variables[0][-6][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-6][1] ) );
    GTECH_OAI2N2 U1143 ( .A(n6350), .B(n6346), .C(\Variables[0][-6][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-6][0] ) );
    GTECH_OAI2N2 U1144 ( .A(n6351), .B(n6346), .C(\Variables[0][-5][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-5][3] ) );
    GTECH_OAI2N2 U1145 ( .A(n6352), .B(n6346), .C(\Variables[0][-5][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-5][2] ) );
    GTECH_OAI2N2 U1146 ( .A(n6353), .B(n6346), .C(\Variables[0][-5][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-5][1] ) );
    GTECH_OAI2N2 U1147 ( .A(n6354), .B(n6346), .C(\Variables[0][-5][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-5][0] ) );
    GTECH_OAI2N2 U1148 ( .A(n6355), .B(n6346), .C(\Variables[0][-4][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-4][3] ) );
    GTECH_OAI2N2 U1149 ( .A(n6356), .B(n6346), .C(\Variables[0][-4][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-4][2] ) );
    GTECH_OAI2N2 U1150 ( .A(n6357), .B(n6346), .C(\Variables[0][-4][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-4][1] ) );
    GTECH_OAI2N2 U1151 ( .A(n6358), .B(n6346), .C(\Variables[0][-4][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-4][0] ) );
    GTECH_NOT U1152 ( .A(n6359), .Z(\Variables2830[0][-3][3] ) );
    GTECH_NOT U1153 ( .A(n6360), .Z(\Variables2830[0][-3][2] ) );
    GTECH_NOT U1154 ( .A(n6361), .Z(\Variables2830[0][-3][1] ) );
    GTECH_NOT U1155 ( .A(n6362), .Z(\Variables2830[0][-3][0] ) );
    GTECH_OAI2N2 U1156 ( .A(n6363), .B(n6346), .C(\Variables[0][-2][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-2][3] ) );
    GTECH_OAI2N2 U1157 ( .A(n6364), .B(n6346), .C(\Variables[0][-2][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-2][2] ) );
    GTECH_OAI2N2 U1158 ( .A(n6365), .B(n6346), .C(\Variables[0][-2][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-2][1] ) );
    GTECH_OAI2N2 U1159 ( .A(n6366), .B(n6346), .C(\Variables[0][-2][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-2][0] ) );
    GTECH_OAI2N2 U1160 ( .A(n6367), .B(n6346), .C(\Variables[0][-1][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-1][3] ) );
    GTECH_OAI2N2 U1161 ( .A(n6368), .B(n6346), .C(\Variables[0][-1][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-1][2] ) );
    GTECH_OAI2N2 U1162 ( .A(n6369), .B(n6346), .C(\Variables[0][-1][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-1][1] ) );
    GTECH_OAI2N2 U1163 ( .A(n6370), .B(n6346), .C(\Variables[0][-1][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][-1][0] ) );
    GTECH_OAI2N2 U1164 ( .A(n6371), .B(n6346), .C(\Variables[0][0][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][0][3] ) );
    GTECH_OAI2N2 U1165 ( .A(n6372), .B(n6346), .C(\Variables[0][0][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][0][2] ) );
    GTECH_OAI2N2 U1166 ( .A(n6373), .B(n6346), .C(\Variables[0][0][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][0][1] ) );
    GTECH_OAI2N2 U1167 ( .A(n6374), .B(n6346), .C(\Variables[0][0][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][0][0] ) );
    GTECH_OAI2N2 U1168 ( .A(n6375), .B(n6346), .C(\Variables[0][1][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][1][3] ) );
    GTECH_OAI2N2 U1169 ( .A(n6376), .B(n6346), .C(\Variables[0][1][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][1][2] ) );
    GTECH_OAI2N2 U1170 ( .A(n6377), .B(n6346), .C(\Variables[0][1][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][1][1] ) );
    GTECH_OAI2N2 U1171 ( .A(n6378), .B(n6346), .C(\Variables[0][1][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][1][0] ) );
    GTECH_OAI2N2 U1172 ( .A(n6379), .B(n6346), .C(\Variables[0][2][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][2][3] ) );
    GTECH_OAI2N2 U1173 ( .A(n6380), .B(n6346), .C(\Variables[0][2][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][2][2] ) );
    GTECH_OAI2N2 U1174 ( .A(n6381), .B(n6346), .C(\Variables[0][2][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][2][1] ) );
    GTECH_OAI2N2 U1175 ( .A(n6382), .B(n6346), .C(\Variables[0][2][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][2][0] ) );
    GTECH_OAI2N2 U1176 ( .A(n6383), .B(n6346), .C(\Variables[0][3][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][3][3] ) );
    GTECH_OAI2N2 U1177 ( .A(n6384), .B(n6346), .C(\Variables[0][3][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][3][2] ) );
    GTECH_OAI2N2 U1178 ( .A(n6385), .B(n6346), .C(\Variables[0][3][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][3][1] ) );
    GTECH_OAI2N2 U1179 ( .A(n6386), .B(n6346), .C(\Variables[0][3][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][3][0] ) );
    GTECH_OAI2N2 U1180 ( .A(n6387), .B(n6346), .C(\Variables[0][4][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][4][3] ) );
    GTECH_OAI2N2 U1181 ( .A(n6388), .B(n6346), .C(\Variables[0][4][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][4][2] ) );
    GTECH_OAI2N2 U1182 ( .A(n6389), .B(n6346), .C(\Variables[0][4][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][4][1] ) );
    GTECH_OAI2N2 U1183 ( .A(n6390), .B(n6346), .C(\Variables[0][4][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][4][0] ) );
    GTECH_OAI2N2 U1184 ( .A(n6391), .B(n6346), .C(\Variables[0][5][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][5][3] ) );
    GTECH_OAI2N2 U1185 ( .A(n6392), .B(n6346), .C(\Variables[0][5][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][5][2] ) );
    GTECH_OAI2N2 U1186 ( .A(n6393), .B(n6346), .C(\Variables[0][5][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][5][1] ) );
    GTECH_OAI2N2 U1187 ( .A(n6394), .B(n6346), .C(\Variables[0][5][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][5][0] ) );
    GTECH_OAI2N2 U1188 ( .A(n6395), .B(n6346), .C(\Variables[0][6][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][6][3] ) );
    GTECH_OAI2N2 U1189 ( .A(n6396), .B(n6346), .C(\Variables[0][6][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][6][2] ) );
    GTECH_OAI2N2 U1190 ( .A(n6397), .B(n6346), .C(\Variables[0][6][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][6][1] ) );
    GTECH_OAI2N2 U1191 ( .A(n6398), .B(n6346), .C(\Variables[0][6][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][6][0] ) );
    GTECH_OAI2N2 U1192 ( .A(n6399), .B(n6346), .C(\Variables[0][7][3]_wire ), 
        .D(n6347), .Z(\Variables2830[0][7][3] ) );
    GTECH_OAI2N2 U1193 ( .A(n6400), .B(n6346), .C(\Variables[0][7][2]_wire ), 
        .D(n6347), .Z(\Variables2830[0][7][2] ) );
    GTECH_OAI2N2 U1194 ( .A(n6401), .B(n6346), .C(\Variables[0][7][1]_wire ), 
        .D(n6347), .Z(\Variables2830[0][7][1] ) );
    GTECH_OAI2N2 U1195 ( .A(n6402), .B(n6346), .C(\Variables[0][7][0]_wire ), 
        .D(n6347), .Z(\Variables2830[0][7][0] ) );
    GTECH_OAI2N2 U1196 ( .A(n6403), .B(n6404), .C(\Variables[1][-8][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-8][3] ) );
    GTECH_OAI2N2 U1197 ( .A(n6406), .B(n6404), .C(\Variables[1][-8][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-8][2] ) );
    GTECH_OAI2N2 U1198 ( .A(n6407), .B(n6404), .C(\Variables[1][-8][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-8][1] ) );
    GTECH_OAI2N2 U1199 ( .A(n6408), .B(n6404), .C(\Variables[1][-8][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-8][0] ) );
    GTECH_OAI2N2 U1200 ( .A(n6409), .B(n6404), .C(\Variables[1][-7][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-7][3] ) );
    GTECH_OAI2N2 U1201 ( .A(n6410), .B(n6404), .C(\Variables[1][-7][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-7][2] ) );
    GTECH_OAI2N2 U1202 ( .A(n6411), .B(n6404), .C(\Variables[1][-7][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-7][1] ) );
    GTECH_OAI2N2 U1203 ( .A(n6412), .B(n6404), .C(\Variables[1][-7][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-7][0] ) );
    GTECH_OAI2N2 U1204 ( .A(n6345), .B(n6404), .C(\Variables[1][-6][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-6][3] ) );
    GTECH_OAI2N2 U1205 ( .A(n6348), .B(n6404), .C(\Variables[1][-6][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-6][2] ) );
    GTECH_OAI2N2 U1206 ( .A(n6349), .B(n6404), .C(\Variables[1][-6][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-6][1] ) );
    GTECH_OAI2N2 U1207 ( .A(n6350), .B(n6404), .C(\Variables[1][-6][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-6][0] ) );
    GTECH_OAI2N2 U1208 ( .A(n6351), .B(n6404), .C(\Variables[1][-5][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-5][3] ) );
    GTECH_OAI2N2 U1209 ( .A(n6352), .B(n6404), .C(\Variables[1][-5][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-5][2] ) );
    GTECH_OAI2N2 U1210 ( .A(n6353), .B(n6404), .C(\Variables[1][-5][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-5][1] ) );
    GTECH_OAI2N2 U1211 ( .A(n6354), .B(n6404), .C(\Variables[1][-5][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-5][0] ) );
    GTECH_OAI2N2 U1212 ( .A(n6355), .B(n6404), .C(\Variables[1][-4][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-4][3] ) );
    GTECH_OAI2N2 U1213 ( .A(n6356), .B(n6404), .C(\Variables[1][-4][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-4][2] ) );
    GTECH_OAI2N2 U1214 ( .A(n6357), .B(n6404), .C(\Variables[1][-4][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-4][1] ) );
    GTECH_OAI2N2 U1215 ( .A(n6358), .B(n6404), .C(\Variables[1][-4][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-4][0] ) );
    GTECH_OAI2N2 U1216 ( .A(n6413), .B(n6404), .C(\Variables[1][-3][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-3][3] ) );
    GTECH_OAI2N2 U1217 ( .A(n6414), .B(n6404), .C(\Variables[1][-3][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-3][2] ) );
    GTECH_OAI2N2 U1218 ( .A(n6415), .B(n6404), .C(\Variables[1][-3][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-3][1] ) );
    GTECH_OAI2N2 U1219 ( .A(n6416), .B(n6404), .C(\Variables[1][-3][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-3][0] ) );
    GTECH_OAI2N2 U1220 ( .A(n6363), .B(n6404), .C(\Variables[1][-2][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-2][3] ) );
    GTECH_OAI2N2 U1221 ( .A(n6364), .B(n6404), .C(\Variables[1][-2][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-2][2] ) );
    GTECH_OAI2N2 U1222 ( .A(n6365), .B(n6404), .C(\Variables[1][-2][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-2][1] ) );
    GTECH_OAI2N2 U1223 ( .A(n6366), .B(n6404), .C(\Variables[1][-2][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-2][0] ) );
    GTECH_OAI2N2 U1224 ( .A(n6367), .B(n6404), .C(\Variables[1][-1][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-1][3] ) );
    GTECH_OAI2N2 U1225 ( .A(n6368), .B(n6404), .C(\Variables[1][-1][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-1][2] ) );
    GTECH_OAI2N2 U1226 ( .A(n6369), .B(n6404), .C(\Variables[1][-1][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-1][1] ) );
    GTECH_OAI2N2 U1227 ( .A(n6370), .B(n6404), .C(\Variables[1][-1][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][-1][0] ) );
    GTECH_OAI2N2 U1228 ( .A(n6371), .B(n6404), .C(\Variables[1][0][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][0][3] ) );
    GTECH_OAI2N2 U1229 ( .A(n6372), .B(n6404), .C(\Variables[1][0][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][0][2] ) );
    GTECH_OAI2N2 U1230 ( .A(n6373), .B(n6404), .C(\Variables[1][0][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][0][1] ) );
    GTECH_OAI2N2 U1231 ( .A(n6374), .B(n6404), .C(\Variables[1][0][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][0][0] ) );
    GTECH_OAI2N2 U1232 ( .A(n6375), .B(n6404), .C(\Variables[1][1][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][1][3] ) );
    GTECH_OAI2N2 U1233 ( .A(n6376), .B(n6404), .C(\Variables[1][1][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][1][2] ) );
    GTECH_OAI2N2 U1234 ( .A(n6377), .B(n6404), .C(\Variables[1][1][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][1][1] ) );
    GTECH_OAI2N2 U1235 ( .A(n6378), .B(n6404), .C(\Variables[1][1][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][1][0] ) );
    GTECH_OAI2N2 U1236 ( .A(n6379), .B(n6404), .C(\Variables[1][2][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][2][3] ) );
    GTECH_OAI2N2 U1237 ( .A(n6380), .B(n6404), .C(\Variables[1][2][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][2][2] ) );
    GTECH_OAI2N2 U1238 ( .A(n6381), .B(n6404), .C(\Variables[1][2][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][2][1] ) );
    GTECH_OAI2N2 U1239 ( .A(n6382), .B(n6404), .C(\Variables[1][2][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][2][0] ) );
    GTECH_OAI2N2 U1240 ( .A(n6383), .B(n6404), .C(\Variables[1][3][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][3][3] ) );
    GTECH_OAI2N2 U1241 ( .A(n6384), .B(n6404), .C(\Variables[1][3][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][3][2] ) );
    GTECH_OAI2N2 U1242 ( .A(n6385), .B(n6404), .C(\Variables[1][3][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][3][1] ) );
    GTECH_OAI2N2 U1243 ( .A(n6386), .B(n6404), .C(\Variables[1][3][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][3][0] ) );
    GTECH_OAI2N2 U1244 ( .A(n6387), .B(n6404), .C(\Variables[1][4][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][4][3] ) );
    GTECH_OAI2N2 U1245 ( .A(n6388), .B(n6404), .C(\Variables[1][4][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][4][2] ) );
    GTECH_OAI2N2 U1246 ( .A(n6389), .B(n6404), .C(\Variables[1][4][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][4][1] ) );
    GTECH_OAI2N2 U1247 ( .A(n6390), .B(n6404), .C(\Variables[1][4][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][4][0] ) );
    GTECH_OAI2N2 U1248 ( .A(n6391), .B(n6404), .C(\Variables[1][5][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][5][3] ) );
    GTECH_OAI2N2 U1249 ( .A(n6392), .B(n6404), .C(\Variables[1][5][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][5][2] ) );
    GTECH_OAI2N2 U1250 ( .A(n6393), .B(n6404), .C(\Variables[1][5][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][5][1] ) );
    GTECH_OAI2N2 U1251 ( .A(n6394), .B(n6404), .C(\Variables[1][5][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][5][0] ) );
    GTECH_OAI2N2 U1252 ( .A(n6395), .B(n6404), .C(\Variables[1][6][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][6][3] ) );
    GTECH_OAI2N2 U1253 ( .A(n6396), .B(n6404), .C(\Variables[1][6][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][6][2] ) );
    GTECH_OAI2N2 U1254 ( .A(n6397), .B(n6404), .C(\Variables[1][6][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][6][1] ) );
    GTECH_OAI2N2 U1255 ( .A(n6398), .B(n6404), .C(\Variables[1][6][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][6][0] ) );
    GTECH_OAI2N2 U1256 ( .A(n6399), .B(n6404), .C(\Variables[1][7][3]_wire ), 
        .D(n6405), .Z(\Variables2830[1][7][3] ) );
    GTECH_OAI2N2 U1257 ( .A(n6400), .B(n6404), .C(\Variables[1][7][2]_wire ), 
        .D(n6405), .Z(\Variables2830[1][7][2] ) );
    GTECH_OAI2N2 U1258 ( .A(n6401), .B(n6404), .C(\Variables[1][7][1]_wire ), 
        .D(n6405), .Z(\Variables2830[1][7][1] ) );
    GTECH_OAI2N2 U1259 ( .A(n6402), .B(n6404), .C(\Variables[1][7][0]_wire ), 
        .D(n6405), .Z(\Variables2830[1][7][0] ) );
    GTECH_OAI2N2 U1260 ( .A(n6403), .B(n6417), .C(\Variables[2][-8][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-8][3] ) );
    GTECH_OAI2N2 U1261 ( .A(n6406), .B(n6417), .C(\Variables[2][-8][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-8][2] ) );
    GTECH_OAI2N2 U1262 ( .A(n6407), .B(n6417), .C(\Variables[2][-8][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-8][1] ) );
    GTECH_OAI2N2 U1263 ( .A(n6408), .B(n6417), .C(\Variables[2][-8][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-8][0] ) );
    GTECH_OAI2N2 U1264 ( .A(n6409), .B(n6417), .C(\Variables[2][-7][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-7][3] ) );
    GTECH_OAI2N2 U1265 ( .A(n6410), .B(n6417), .C(\Variables[2][-7][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-7][2] ) );
    GTECH_OAI2N2 U1266 ( .A(n6411), .B(n6417), .C(\Variables[2][-7][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-7][1] ) );
    GTECH_OAI2N2 U1267 ( .A(n6412), .B(n6417), .C(\Variables[2][-7][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-7][0] ) );
    GTECH_OAI2N2 U1268 ( .A(n6345), .B(n6417), .C(\Variables[2][-6][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-6][3] ) );
    GTECH_OAI2N2 U1269 ( .A(n6348), .B(n6417), .C(\Variables[2][-6][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-6][2] ) );
    GTECH_OAI2N2 U1270 ( .A(n6349), .B(n6417), .C(\Variables[2][-6][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-6][1] ) );
    GTECH_OAI2N2 U1271 ( .A(n6350), .B(n6417), .C(\Variables[2][-6][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-6][0] ) );
    GTECH_OAI2N2 U1272 ( .A(n6351), .B(n6417), .C(\Variables[2][-5][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-5][3] ) );
    GTECH_OAI2N2 U1273 ( .A(n6352), .B(n6417), .C(\Variables[2][-5][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-5][2] ) );
    GTECH_OAI2N2 U1274 ( .A(n6353), .B(n6417), .C(\Variables[2][-5][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-5][1] ) );
    GTECH_OAI2N2 U1275 ( .A(n6354), .B(n6417), .C(\Variables[2][-5][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-5][0] ) );
    GTECH_OAI2N2 U1276 ( .A(n6355), .B(n6417), .C(\Variables[2][-4][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-4][3] ) );
    GTECH_OAI2N2 U1277 ( .A(n6356), .B(n6417), .C(\Variables[2][-4][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-4][2] ) );
    GTECH_OAI2N2 U1278 ( .A(n6357), .B(n6417), .C(\Variables[2][-4][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-4][1] ) );
    GTECH_OAI2N2 U1279 ( .A(n6358), .B(n6417), .C(\Variables[2][-4][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-4][0] ) );
    GTECH_OAI2N2 U1280 ( .A(n6413), .B(n6417), .C(\Variables[2][-3][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-3][3] ) );
    GTECH_OAI2N2 U1281 ( .A(n6414), .B(n6417), .C(\Variables[2][-3][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-3][2] ) );
    GTECH_OAI2N2 U1282 ( .A(n6415), .B(n6417), .C(\Variables[2][-3][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-3][1] ) );
    GTECH_OAI2N2 U1283 ( .A(n6416), .B(n6417), .C(\Variables[2][-3][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-3][0] ) );
    GTECH_OAI2N2 U1284 ( .A(n6363), .B(n6417), .C(\Variables[2][-2][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-2][3] ) );
    GTECH_OAI2N2 U1285 ( .A(n6364), .B(n6417), .C(\Variables[2][-2][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-2][2] ) );
    GTECH_OAI2N2 U1286 ( .A(n6365), .B(n6417), .C(\Variables[2][-2][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-2][1] ) );
    GTECH_OAI2N2 U1287 ( .A(n6366), .B(n6417), .C(\Variables[2][-2][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-2][0] ) );
    GTECH_OAI2N2 U1288 ( .A(n6367), .B(n6417), .C(\Variables[2][-1][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-1][3] ) );
    GTECH_OAI2N2 U1289 ( .A(n6368), .B(n6417), .C(\Variables[2][-1][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-1][2] ) );
    GTECH_OAI2N2 U1290 ( .A(n6369), .B(n6417), .C(\Variables[2][-1][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-1][1] ) );
    GTECH_OAI2N2 U1291 ( .A(n6370), .B(n6417), .C(\Variables[2][-1][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][-1][0] ) );
    GTECH_OAI2N2 U1292 ( .A(n6371), .B(n6417), .C(\Variables[2][0][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][0][3] ) );
    GTECH_OAI2N2 U1293 ( .A(n6372), .B(n6417), .C(\Variables[2][0][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][0][2] ) );
    GTECH_OAI2N2 U1294 ( .A(n6373), .B(n6417), .C(\Variables[2][0][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][0][1] ) );
    GTECH_OAI2N2 U1295 ( .A(n6374), .B(n6417), .C(\Variables[2][0][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][0][0] ) );
    GTECH_OAI2N2 U1296 ( .A(n6375), .B(n6417), .C(\Variables[2][1][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][1][3] ) );
    GTECH_OAI2N2 U1297 ( .A(n6376), .B(n6417), .C(\Variables[2][1][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][1][2] ) );
    GTECH_OAI2N2 U1298 ( .A(n6377), .B(n6417), .C(\Variables[2][1][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][1][1] ) );
    GTECH_OAI2N2 U1299 ( .A(n6378), .B(n6417), .C(\Variables[2][1][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][1][0] ) );
    GTECH_OAI2N2 U1300 ( .A(n6379), .B(n6417), .C(\Variables[2][2][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][2][3] ) );
    GTECH_OAI2N2 U1301 ( .A(n6380), .B(n6417), .C(\Variables[2][2][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][2][2] ) );
    GTECH_OAI2N2 U1302 ( .A(n6381), .B(n6417), .C(\Variables[2][2][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][2][1] ) );
    GTECH_OAI2N2 U1303 ( .A(n6382), .B(n6417), .C(\Variables[2][2][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][2][0] ) );
    GTECH_OAI2N2 U1304 ( .A(n6383), .B(n6417), .C(\Variables[2][3][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][3][3] ) );
    GTECH_OAI2N2 U1305 ( .A(n6384), .B(n6417), .C(\Variables[2][3][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][3][2] ) );
    GTECH_OAI2N2 U1306 ( .A(n6385), .B(n6417), .C(\Variables[2][3][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][3][1] ) );
    GTECH_OAI2N2 U1307 ( .A(n6386), .B(n6417), .C(\Variables[2][3][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][3][0] ) );
    GTECH_OAI2N2 U1308 ( .A(n6387), .B(n6417), .C(\Variables[2][4][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][4][3] ) );
    GTECH_OAI2N2 U1309 ( .A(n6388), .B(n6417), .C(\Variables[2][4][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][4][2] ) );
    GTECH_OAI2N2 U1310 ( .A(n6389), .B(n6417), .C(\Variables[2][4][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][4][1] ) );
    GTECH_OAI2N2 U1311 ( .A(n6390), .B(n6417), .C(\Variables[2][4][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][4][0] ) );
    GTECH_OAI2N2 U1312 ( .A(n6391), .B(n6417), .C(\Variables[2][5][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][5][3] ) );
    GTECH_OAI2N2 U1313 ( .A(n6392), .B(n6417), .C(\Variables[2][5][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][5][2] ) );
    GTECH_OAI2N2 U1314 ( .A(n6393), .B(n6417), .C(\Variables[2][5][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][5][1] ) );
    GTECH_OAI2N2 U1315 ( .A(n6394), .B(n6417), .C(\Variables[2][5][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][5][0] ) );
    GTECH_OAI2N2 U1316 ( .A(n6395), .B(n6417), .C(\Variables[2][6][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][6][3] ) );
    GTECH_OAI2N2 U1317 ( .A(n6396), .B(n6417), .C(\Variables[2][6][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][6][2] ) );
    GTECH_OAI2N2 U1318 ( .A(n6397), .B(n6417), .C(\Variables[2][6][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][6][1] ) );
    GTECH_OAI2N2 U1319 ( .A(n6398), .B(n6417), .C(\Variables[2][6][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][6][0] ) );
    GTECH_OAI2N2 U1320 ( .A(n6399), .B(n6417), .C(\Variables[2][7][3]_wire ), 
        .D(n6418), .Z(\Variables2830[2][7][3] ) );
    GTECH_OAI2N2 U1321 ( .A(n6400), .B(n6417), .C(\Variables[2][7][2]_wire ), 
        .D(n6418), .Z(\Variables2830[2][7][2] ) );
    GTECH_OAI2N2 U1322 ( .A(n6401), .B(n6417), .C(\Variables[2][7][1]_wire ), 
        .D(n6418), .Z(\Variables2830[2][7][1] ) );
    GTECH_OAI2N2 U1323 ( .A(n6402), .B(n6417), .C(\Variables[2][7][0]_wire ), 
        .D(n6418), .Z(\Variables2830[2][7][0] ) );
    GTECH_OAI2N2 U1324 ( .A(n6403), .B(n6419), .C(\Variables[3][-8][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-8][3] ) );
    GTECH_OAI2N2 U1325 ( .A(n6406), .B(n6419), .C(\Variables[3][-8][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-8][2] ) );
    GTECH_OAI2N2 U1326 ( .A(n6407), .B(n6419), .C(\Variables[3][-8][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-8][1] ) );
    GTECH_OAI2N2 U1327 ( .A(n6408), .B(n6419), .C(\Variables[3][-8][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-8][0] ) );
    GTECH_OAI2N2 U1328 ( .A(n6409), .B(n6419), .C(\Variables[3][-7][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-7][3] ) );
    GTECH_OAI2N2 U1329 ( .A(n6410), .B(n6419), .C(\Variables[3][-7][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-7][2] ) );
    GTECH_OAI2N2 U1330 ( .A(n6411), .B(n6419), .C(\Variables[3][-7][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-7][1] ) );
    GTECH_OAI2N2 U1331 ( .A(n6412), .B(n6419), .C(\Variables[3][-7][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-7][0] ) );
    GTECH_OAI2N2 U1332 ( .A(n6345), .B(n6419), .C(\Variables[3][-6][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-6][3] ) );
    GTECH_OAI2N2 U1333 ( .A(n6348), .B(n6419), .C(\Variables[3][-6][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-6][2] ) );
    GTECH_OAI2N2 U1334 ( .A(n6349), .B(n6419), .C(\Variables[3][-6][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-6][1] ) );
    GTECH_OAI2N2 U1335 ( .A(n6350), .B(n6419), .C(\Variables[3][-6][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-6][0] ) );
    GTECH_OAI2N2 U1336 ( .A(n6351), .B(n6419), .C(\Variables[3][-5][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-5][3] ) );
    GTECH_OAI2N2 U1337 ( .A(n6352), .B(n6419), .C(\Variables[3][-5][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-5][2] ) );
    GTECH_OAI2N2 U1338 ( .A(n6353), .B(n6419), .C(\Variables[3][-5][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-5][1] ) );
    GTECH_OAI2N2 U1339 ( .A(n6354), .B(n6419), .C(\Variables[3][-5][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-5][0] ) );
    GTECH_OAI2N2 U1340 ( .A(n6355), .B(n6419), .C(\Variables[3][-4][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-4][3] ) );
    GTECH_OAI2N2 U1341 ( .A(n6356), .B(n6419), .C(\Variables[3][-4][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-4][2] ) );
    GTECH_OAI2N2 U1342 ( .A(n6357), .B(n6419), .C(\Variables[3][-4][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-4][1] ) );
    GTECH_OAI2N2 U1343 ( .A(n6358), .B(n6419), .C(\Variables[3][-4][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-4][0] ) );
    GTECH_OAI2N2 U1344 ( .A(n6413), .B(n6419), .C(\Variables[3][-3][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-3][3] ) );
    GTECH_OAI2N2 U1345 ( .A(n6414), .B(n6419), .C(\Variables[3][-3][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-3][2] ) );
    GTECH_OAI2N2 U1346 ( .A(n6415), .B(n6419), .C(\Variables[3][-3][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-3][1] ) );
    GTECH_OAI2N2 U1347 ( .A(n6416), .B(n6419), .C(\Variables[3][-3][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-3][0] ) );
    GTECH_OAI2N2 U1348 ( .A(n6363), .B(n6419), .C(\Variables[3][-2][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-2][3] ) );
    GTECH_OAI2N2 U1349 ( .A(n6364), .B(n6419), .C(\Variables[3][-2][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-2][2] ) );
    GTECH_OAI2N2 U1350 ( .A(n6365), .B(n6419), .C(\Variables[3][-2][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-2][1] ) );
    GTECH_OAI2N2 U1351 ( .A(n6366), .B(n6419), .C(\Variables[3][-2][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-2][0] ) );
    GTECH_OAI2N2 U1352 ( .A(n6367), .B(n6419), .C(\Variables[3][-1][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-1][3] ) );
    GTECH_OAI2N2 U1353 ( .A(n6368), .B(n6419), .C(\Variables[3][-1][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-1][2] ) );
    GTECH_OAI2N2 U1354 ( .A(n6369), .B(n6419), .C(\Variables[3][-1][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-1][1] ) );
    GTECH_OAI2N2 U1355 ( .A(n6370), .B(n6419), .C(\Variables[3][-1][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][-1][0] ) );
    GTECH_OAI2N2 U1356 ( .A(n6371), .B(n6419), .C(\Variables[3][0][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][0][3] ) );
    GTECH_OAI2N2 U1357 ( .A(n6372), .B(n6419), .C(\Variables[3][0][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][0][2] ) );
    GTECH_OAI2N2 U1358 ( .A(n6373), .B(n6419), .C(\Variables[3][0][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][0][1] ) );
    GTECH_OAI2N2 U1359 ( .A(n6374), .B(n6419), .C(\Variables[3][0][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][0][0] ) );
    GTECH_OAI2N2 U1360 ( .A(n6375), .B(n6419), .C(\Variables[3][1][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][1][3] ) );
    GTECH_OAI2N2 U1361 ( .A(n6376), .B(n6419), .C(\Variables[3][1][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][1][2] ) );
    GTECH_OAI2N2 U1362 ( .A(n6377), .B(n6419), .C(\Variables[3][1][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][1][1] ) );
    GTECH_OAI2N2 U1363 ( .A(n6378), .B(n6419), .C(\Variables[3][1][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][1][0] ) );
    GTECH_OAI2N2 U1364 ( .A(n6379), .B(n6419), .C(\Variables[3][2][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][2][3] ) );
    GTECH_OAI2N2 U1365 ( .A(n6380), .B(n6419), .C(\Variables[3][2][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][2][2] ) );
    GTECH_OAI2N2 U1366 ( .A(n6381), .B(n6419), .C(\Variables[3][2][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][2][1] ) );
    GTECH_OAI2N2 U1367 ( .A(n6382), .B(n6419), .C(\Variables[3][2][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][2][0] ) );
    GTECH_OAI2N2 U1368 ( .A(n6383), .B(n6419), .C(\Variables[3][3][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][3][3] ) );
    GTECH_OAI2N2 U1369 ( .A(n6384), .B(n6419), .C(\Variables[3][3][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][3][2] ) );
    GTECH_OAI2N2 U1370 ( .A(n6385), .B(n6419), .C(\Variables[3][3][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][3][1] ) );
    GTECH_OAI2N2 U1371 ( .A(n6386), .B(n6419), .C(\Variables[3][3][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][3][0] ) );
    GTECH_OAI2N2 U1372 ( .A(n6387), .B(n6419), .C(\Variables[3][4][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][4][3] ) );
    GTECH_OAI2N2 U1373 ( .A(n6388), .B(n6419), .C(\Variables[3][4][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][4][2] ) );
    GTECH_OAI2N2 U1374 ( .A(n6389), .B(n6419), .C(\Variables[3][4][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][4][1] ) );
    GTECH_OAI2N2 U1375 ( .A(n6390), .B(n6419), .C(\Variables[3][4][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][4][0] ) );
    GTECH_OAI2N2 U1376 ( .A(n6391), .B(n6419), .C(\Variables[3][5][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][5][3] ) );
    GTECH_OAI2N2 U1377 ( .A(n6392), .B(n6419), .C(\Variables[3][5][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][5][2] ) );
    GTECH_OAI2N2 U1378 ( .A(n6393), .B(n6419), .C(\Variables[3][5][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][5][1] ) );
    GTECH_OAI2N2 U1379 ( .A(n6394), .B(n6419), .C(\Variables[3][5][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][5][0] ) );
    GTECH_OAI2N2 U1380 ( .A(n6395), .B(n6419), .C(\Variables[3][6][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][6][3] ) );
    GTECH_OAI2N2 U1381 ( .A(n6396), .B(n6419), .C(\Variables[3][6][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][6][2] ) );
    GTECH_OAI2N2 U1382 ( .A(n6397), .B(n6419), .C(\Variables[3][6][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][6][1] ) );
    GTECH_OAI2N2 U1383 ( .A(n6398), .B(n6419), .C(\Variables[3][6][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][6][0] ) );
    GTECH_OAI2N2 U1384 ( .A(n6399), .B(n6419), .C(\Variables[3][7][3]_wire ), 
        .D(n6420), .Z(\Variables2830[3][7][3] ) );
    GTECH_OAI2N2 U1385 ( .A(n6400), .B(n6419), .C(\Variables[3][7][2]_wire ), 
        .D(n6420), .Z(\Variables2830[3][7][2] ) );
    GTECH_OAI2N2 U1386 ( .A(n6401), .B(n6419), .C(\Variables[3][7][1]_wire ), 
        .D(n6420), .Z(\Variables2830[3][7][1] ) );
    GTECH_OAI2N2 U1387 ( .A(n6402), .B(n6419), .C(\Variables[3][7][0]_wire ), 
        .D(n6420), .Z(\Variables2830[3][7][0] ) );
    GTECH_OAI2N2 U1388 ( .A(n6403), .B(n6421), .C(n6422), .D(
        \Variables[4][-8][3]_wire ), .Z(\Variables2830[4][-8][3] ) );
    GTECH_OAI2N2 U1389 ( .A(n6406), .B(n6421), .C(n6422), .D(
        \Variables[4][-8][2]_wire ), .Z(\Variables2830[4][-8][2] ) );
    GTECH_OAI2N2 U1390 ( .A(n6407), .B(n6421), .C(n6422), .D(
        \Variables[4][-8][1]_wire ), .Z(\Variables2830[4][-8][1] ) );
    GTECH_OAI2N2 U1391 ( .A(n6408), .B(n6421), .C(n6422), .D(
        \Variables[4][-8][0]_wire ), .Z(\Variables2830[4][-8][0] ) );
    GTECH_OAI2N2 U1392 ( .A(n6409), .B(n6421), .C(n6422), .D(
        \Variables[4][-7][3]_wire ), .Z(\Variables2830[4][-7][3] ) );
    GTECH_OAI2N2 U1393 ( .A(n6410), .B(n6421), .C(n6422), .D(
        \Variables[4][-7][2]_wire ), .Z(\Variables2830[4][-7][2] ) );
    GTECH_OAI2N2 U1394 ( .A(n6411), .B(n6421), .C(n6422), .D(
        \Variables[4][-7][1]_wire ), .Z(\Variables2830[4][-7][1] ) );
    GTECH_OAI2N2 U1395 ( .A(n6412), .B(n6421), .C(n6422), .D(
        \Variables[4][-7][0]_wire ), .Z(\Variables2830[4][-7][0] ) );
    GTECH_OAI2N2 U1396 ( .A(n6345), .B(n6421), .C(n6422), .D(
        \Variables[4][-6][3]_wire ), .Z(\Variables2830[4][-6][3] ) );
    GTECH_OAI2N2 U1397 ( .A(n6348), .B(n6421), .C(n6422), .D(
        \Variables[4][-6][2]_wire ), .Z(\Variables2830[4][-6][2] ) );
    GTECH_OAI2N2 U1398 ( .A(n6349), .B(n6421), .C(n6422), .D(
        \Variables[4][-6][1]_wire ), .Z(\Variables2830[4][-6][1] ) );
    GTECH_OAI2N2 U1399 ( .A(n6350), .B(n6421), .C(n6422), .D(
        \Variables[4][-6][0]_wire ), .Z(\Variables2830[4][-6][0] ) );
    GTECH_OAI2N2 U1400 ( .A(n6351), .B(n6421), .C(n6422), .D(
        \Variables[4][-5][3]_wire ), .Z(\Variables2830[4][-5][3] ) );
    GTECH_OAI2N2 U1401 ( .A(n6352), .B(n6421), .C(n6422), .D(
        \Variables[4][-5][2]_wire ), .Z(\Variables2830[4][-5][2] ) );
    GTECH_OAI2N2 U1402 ( .A(n6353), .B(n6421), .C(n6422), .D(
        \Variables[4][-5][1]_wire ), .Z(\Variables2830[4][-5][1] ) );
    GTECH_OAI2N2 U1403 ( .A(n6354), .B(n6421), .C(n6422), .D(
        \Variables[4][-5][0]_wire ), .Z(\Variables2830[4][-5][0] ) );
    GTECH_OAI2N2 U1404 ( .A(n6355), .B(n6421), .C(n6422), .D(
        \Variables[4][-4][3]_wire ), .Z(\Variables2830[4][-4][3] ) );
    GTECH_OAI2N2 U1405 ( .A(n6356), .B(n6421), .C(n6422), .D(
        \Variables[4][-4][2]_wire ), .Z(\Variables2830[4][-4][2] ) );
    GTECH_OAI2N2 U1406 ( .A(n6357), .B(n6421), .C(n6422), .D(
        \Variables[4][-4][1]_wire ), .Z(\Variables2830[4][-4][1] ) );
    GTECH_OAI2N2 U1407 ( .A(n6358), .B(n6421), .C(n6422), .D(
        \Variables[4][-4][0]_wire ), .Z(\Variables2830[4][-4][0] ) );
    GTECH_OAI2N2 U1408 ( .A(n6413), .B(n6421), .C(n6422), .D(
        \Variables[4][-3][3]_wire ), .Z(\Variables2830[4][-3][3] ) );
    GTECH_OAI2N2 U1409 ( .A(n6414), .B(n6421), .C(n6422), .D(
        \Variables[4][-3][2]_wire ), .Z(\Variables2830[4][-3][2] ) );
    GTECH_OAI2N2 U1410 ( .A(n6415), .B(n6421), .C(n6422), .D(
        \Variables[4][-3][1]_wire ), .Z(\Variables2830[4][-3][1] ) );
    GTECH_OAI2N2 U1411 ( .A(n6416), .B(n6421), .C(n6422), .D(
        \Variables[4][-3][0]_wire ), .Z(\Variables2830[4][-3][0] ) );
    GTECH_OAI2N2 U1412 ( .A(n6363), .B(n6421), .C(n6422), .D(
        \Variables[4][-2][3]_wire ), .Z(\Variables2830[4][-2][3] ) );
    GTECH_OAI2N2 U1413 ( .A(n6364), .B(n6421), .C(n6422), .D(
        \Variables[4][-2][2]_wire ), .Z(\Variables2830[4][-2][2] ) );
    GTECH_OAI2N2 U1414 ( .A(n6365), .B(n6421), .C(n6422), .D(
        \Variables[4][-2][1]_wire ), .Z(\Variables2830[4][-2][1] ) );
    GTECH_OAI2N2 U1415 ( .A(n6366), .B(n6421), .C(n6422), .D(
        \Variables[4][-2][0]_wire ), .Z(\Variables2830[4][-2][0] ) );
    GTECH_OAI2N2 U1416 ( .A(n6367), .B(n6421), .C(n6422), .D(
        \Variables[4][-1][3]_wire ), .Z(\Variables2830[4][-1][3] ) );
    GTECH_OAI2N2 U1417 ( .A(n6368), .B(n6421), .C(n6422), .D(
        \Variables[4][-1][2]_wire ), .Z(\Variables2830[4][-1][2] ) );
    GTECH_OAI2N2 U1418 ( .A(n6369), .B(n6421), .C(n6422), .D(
        \Variables[4][-1][1]_wire ), .Z(\Variables2830[4][-1][1] ) );
    GTECH_OAI2N2 U1419 ( .A(n6370), .B(n6421), .C(n6422), .D(
        \Variables[4][-1][0]_wire ), .Z(\Variables2830[4][-1][0] ) );
    GTECH_OAI2N2 U1420 ( .A(n6371), .B(n6421), .C(n6422), .D(
        \Variables[4][0][3]_wire ), .Z(\Variables2830[4][0][3] ) );
    GTECH_OAI2N2 U1421 ( .A(n6372), .B(n6421), .C(n6422), .D(
        \Variables[4][0][2]_wire ), .Z(\Variables2830[4][0][2] ) );
    GTECH_OAI2N2 U1422 ( .A(n6373), .B(n6421), .C(n6422), .D(
        \Variables[4][0][1]_wire ), .Z(\Variables2830[4][0][1] ) );
    GTECH_OAI2N2 U1423 ( .A(n6374), .B(n6421), .C(n6422), .D(
        \Variables[4][0][0]_wire ), .Z(\Variables2830[4][0][0] ) );
    GTECH_OAI2N2 U1424 ( .A(n6375), .B(n6421), .C(n6422), .D(
        \Variables[4][1][3]_wire ), .Z(\Variables2830[4][1][3] ) );
    GTECH_OAI2N2 U1425 ( .A(n6376), .B(n6421), .C(n6422), .D(
        \Variables[4][1][2]_wire ), .Z(\Variables2830[4][1][2] ) );
    GTECH_OAI2N2 U1426 ( .A(n6377), .B(n6421), .C(n6422), .D(
        \Variables[4][1][1]_wire ), .Z(\Variables2830[4][1][1] ) );
    GTECH_OAI2N2 U1427 ( .A(n6378), .B(n6421), .C(n6422), .D(
        \Variables[4][1][0]_wire ), .Z(\Variables2830[4][1][0] ) );
    GTECH_OAI2N2 U1428 ( .A(n6379), .B(n6421), .C(n6422), .D(
        \Variables[4][2][3]_wire ), .Z(\Variables2830[4][2][3] ) );
    GTECH_OAI2N2 U1429 ( .A(n6380), .B(n6421), .C(n6422), .D(
        \Variables[4][2][2]_wire ), .Z(\Variables2830[4][2][2] ) );
    GTECH_OAI2N2 U1430 ( .A(n6381), .B(n6421), .C(n6422), .D(
        \Variables[4][2][1]_wire ), .Z(\Variables2830[4][2][1] ) );
    GTECH_OAI2N2 U1431 ( .A(n6382), .B(n6421), .C(n6422), .D(
        \Variables[4][2][0]_wire ), .Z(\Variables2830[4][2][0] ) );
    GTECH_OAI2N2 U1432 ( .A(n6383), .B(n6421), .C(n6422), .D(
        \Variables[4][3][3]_wire ), .Z(\Variables2830[4][3][3] ) );
    GTECH_OAI2N2 U1433 ( .A(n6384), .B(n6421), .C(n6422), .D(
        \Variables[4][3][2]_wire ), .Z(\Variables2830[4][3][2] ) );
    GTECH_OAI2N2 U1434 ( .A(n6385), .B(n6421), .C(n6422), .D(
        \Variables[4][3][1]_wire ), .Z(\Variables2830[4][3][1] ) );
    GTECH_OAI2N2 U1435 ( .A(n6386), .B(n6421), .C(n6422), .D(
        \Variables[4][3][0]_wire ), .Z(\Variables2830[4][3][0] ) );
    GTECH_OAI2N2 U1436 ( .A(n6387), .B(n6421), .C(n6422), .D(
        \Variables[4][4][3]_wire ), .Z(\Variables2830[4][4][3] ) );
    GTECH_OAI2N2 U1437 ( .A(n6388), .B(n6421), .C(n6422), .D(
        \Variables[4][4][2]_wire ), .Z(\Variables2830[4][4][2] ) );
    GTECH_OAI2N2 U1438 ( .A(n6389), .B(n6421), .C(n6422), .D(
        \Variables[4][4][1]_wire ), .Z(\Variables2830[4][4][1] ) );
    GTECH_OAI2N2 U1439 ( .A(n6390), .B(n6421), .C(n6422), .D(
        \Variables[4][4][0]_wire ), .Z(\Variables2830[4][4][0] ) );
    GTECH_OAI2N2 U1440 ( .A(n6391), .B(n6421), .C(n6422), .D(
        \Variables[4][5][3]_wire ), .Z(\Variables2830[4][5][3] ) );
    GTECH_OAI2N2 U1441 ( .A(n6392), .B(n6421), .C(n6422), .D(
        \Variables[4][5][2]_wire ), .Z(\Variables2830[4][5][2] ) );
    GTECH_OAI2N2 U1442 ( .A(n6393), .B(n6421), .C(n6422), .D(
        \Variables[4][5][1]_wire ), .Z(\Variables2830[4][5][1] ) );
    GTECH_OAI2N2 U1443 ( .A(n6394), .B(n6421), .C(n6422), .D(
        \Variables[4][5][0]_wire ), .Z(\Variables2830[4][5][0] ) );
    GTECH_OAI2N2 U1444 ( .A(n6395), .B(n6421), .C(n6422), .D(
        \Variables[4][6][3]_wire ), .Z(\Variables2830[4][6][3] ) );
    GTECH_OAI2N2 U1445 ( .A(n6396), .B(n6421), .C(n6422), .D(
        \Variables[4][6][2]_wire ), .Z(\Variables2830[4][6][2] ) );
    GTECH_OAI2N2 U1446 ( .A(n6397), .B(n6421), .C(n6422), .D(
        \Variables[4][6][1]_wire ), .Z(\Variables2830[4][6][1] ) );
    GTECH_OAI2N2 U1447 ( .A(n6398), .B(n6421), .C(n6422), .D(
        \Variables[4][6][0]_wire ), .Z(\Variables2830[4][6][0] ) );
    GTECH_OAI2N2 U1448 ( .A(n6399), .B(n6421), .C(n6422), .D(
        \Variables[4][7][3]_wire ), .Z(\Variables2830[4][7][3] ) );
    GTECH_OAI2N2 U1449 ( .A(n6400), .B(n6421), .C(n6422), .D(
        \Variables[4][7][2]_wire ), .Z(\Variables2830[4][7][2] ) );
    GTECH_OAI2N2 U1450 ( .A(n6401), .B(n6421), .C(n6422), .D(
        \Variables[4][7][1]_wire ), .Z(\Variables2830[4][7][1] ) );
    GTECH_OAI2N2 U1451 ( .A(n6402), .B(n6421), .C(n6422), .D(
        \Variables[4][7][0]_wire ), .Z(\Variables2830[4][7][0] ) );
    GTECH_NAND2 U1452 ( .A(n6423), .B(n6424), .Z(\n2831[0][-8][3] ) );
    GTECH_NAND2 U1453 ( .A(n6423), .B(n6425), .Z(\n2831[0][-3][3] ) );
    GTECH_OAI21 U1454 ( .A(ResetStarted), .B(n6331), .C(n6426), .Z(
        IRQInProcess602) );
    GTECH_OAI21 U1455 ( .A(n6427), .B(n6428), .C(n6429), .Z(n603) );
    GTECH_AND2 U1456 ( .A(n6430), .B(n6431), .Z(IRQWait611) );
    GTECH_OAI21 U1457 ( .A(n6432), .B(n6428), .C(n6429), .Z(n612) );
    GTECH_AND2 U1458 ( .A(\sum1105[2] ), .B(n6322), .Z(\ClockCycleCount621[2] 
        ) );
    GTECH_AND2 U1459 ( .A(\sum1105[1] ), .B(n6322), .Z(\ClockCycleCount621[1] 
        ) );
    GTECH_OAI2N2 U1460 ( .A(n6433), .B(n6434), .C(MemoryReadValue[7]), .D(
        n6435), .Z(\Answer2629[3] ) );
    GTECH_OAI2N2 U1461 ( .A(n6436), .B(n6434), .C(MemoryReadValue[6]), .D(
        n6435), .Z(\Answer2629[2] ) );
    GTECH_OAI2N2 U1462 ( .A(n6437), .B(n6434), .C(MemoryReadValue[5]), .D(
        n6435), .Z(\Answer2629[1] ) );
    GTECH_OAI2N2 U1463 ( .A(n6438), .B(n6434), .C(MemoryReadValue[4]), .D(
        n6435), .Z(\Answer2629[0] ) );
    GTECH_AO21 U1464 ( .A(MemoryReady), .B(Read_wire), .C(n6439), .Z(\n630[3] 
        ) );
    GTECH_OAI21 U1465 ( .A(n6426), .B(n6440), .C(n6441), .Z(\Answer639[3] ) );
    GTECH_OAI21 U1466 ( .A(n6426), .B(n6442), .C(n6443), .Z(\Answer639[2] ) );
    GTECH_OAI21 U1467 ( .A(n6426), .B(n6444), .C(n6445), .Z(\Answer639[1] ) );
    GTECH_OAI21 U1468 ( .A(n6426), .B(n6446), .C(n6447), .Z(\Answer639[0] ) );
    GTECH_AND2 U1469 ( .A(n6430), .B(n6448), .Z(Read648) );
    GTECH_AND2 U1470 ( .A(n6430), .B(n6449), .Z(Write657) );
    GTECH_OAI21 U1471 ( .A(n6450), .B(n6451), .C(n6452), .Z(
        \TableSelect667[3] ) );
    GTECH_OAI21 U1472 ( .A(n6453), .B(n6451), .C(n6454), .Z(
        \TableSelect667[2] ) );
    GTECH_OAI22 U1473 ( .A(\NextInstruction[INSTRUCTION][1] ), .B(
        IRQCLKEnable676), .C(n6455), .D(n6451), .Z(\TableSelect667[1] ) );
    GTECH_OAI22 U1474 ( .A(\NextInstruction[INSTRUCTION][1] ), .B(IRQEnable685
        ), .C(n6456), .D(n6451), .Z(\TableSelect667[0] ) );
    GTECH_NAND3 U1475 ( .A(n6457), .B(n6322), .C(n6458), .Z(\n668[3] ) );
    GTECH_NAND2 U1476 ( .A(\NextInstruction[PARAMETER][1] ), .B(n6322), .Z(
        IRQCLKEnable676) );
    GTECH_NAND2 U1477 ( .A(n6322), .B(n6459), .Z(n677) );
    GTECH_NAND2 U1478 ( .A(\NextInstruction[PARAMETER][0] ), .B(n6322), .Z(
        IRQEnable685) );
    GTECH_AO21 U1479 ( .A(n6329), .B(n6460), .C(ResetStarted), .Z(n686) );
    GTECH_AND2 U1480 ( .A(\*cell*469/U7/Z_0 ), .B(n6322), .Z(\n696[3] ) );
    GTECH_AND2 U1481 ( .A(\*cell*469/U12/Z_0 ), .B(n6322), .Z(\n706[3] ) );
    GTECH_OR3 U1482 ( .A(MemoryReady), .B(ResetStarted), .C(\n3651[7] ), .Z(
        n3641) );
    GTECH_OR_NOT U1483 ( .A(n_324), .B(n7346), .Z(\*cell*469/U144/Z_0 ) );
    GTECH_NOT U1484 ( .A(n_324), .Z(n_323) );
    GTECH_OAI2N2 U1485 ( .A(n6461), .B(n6462), .C(n6463), .D(\sum2964[7] ), 
        .Z(\InstructionPtr3995[7] ) );
    GTECH_OAI2N2 U1486 ( .A(n6464), .B(n6462), .C(n6463), .D(\sum2964[6] ), 
        .Z(\InstructionPtr3995[6] ) );
    GTECH_OAI2N2 U1487 ( .A(n6465), .B(n6462), .C(n6463), .D(\sum2964[5] ), 
        .Z(\InstructionPtr3995[5] ) );
    GTECH_OAI2N2 U1488 ( .A(n6466), .B(n6462), .C(n6463), .D(\sum2964[4] ), 
        .Z(\InstructionPtr3995[4] ) );
    GTECH_OAI2N2 U1489 ( .A(n6467), .B(n6462), .C(n6463), .D(\sum2964[3] ), 
        .Z(\InstructionPtr3995[3] ) );
    GTECH_OAI2N2 U1490 ( .A(n6468), .B(n6462), .C(n6463), .D(\sum2964[2] ), 
        .Z(\InstructionPtr3995[2] ) );
    GTECH_OAI2N2 U1491 ( .A(n6469), .B(n6462), .C(n6463), .D(\sum2964[1] ), 
        .Z(\InstructionPtr3995[1] ) );
    GTECH_OAI2N2 U1492 ( .A(n6470), .B(n6462), .C(n6463), .D(\sum2964[0] ), 
        .Z(\InstructionPtr3995[0] ) );
    GTECH_NAND2 U1493 ( .A(n6471), .B(n6463), .Z(\n3996[7] ) );
    GTECH_OR_NOT U1494 ( .A(n_168), .B(n7335), .Z(\CycleWaveform34[5] ) );
    GTECH_OAI21 U1495 ( .A(ResetStarted), .B(n7330), .C(n6472), .Z(
        \CycleWaveform34[4] ) );
    GTECH_OAI21 U1496 ( .A(ResetStarted), .B(n7331), .C(n6472), .Z(
        \CycleWaveform34[3] ) );
    GTECH_OAI21 U1497 ( .A(ResetStarted), .B(n7332), .C(n6472), .Z(
        \CycleWaveform34[2] ) );
    GTECH_OAI21 U1498 ( .A(ResetStarted), .B(n7333), .C(n6472), .Z(
        \CycleWaveform34[1] ) );
    GTECH_OAI21 U1499 ( .A(ResetStarted), .B(n7334), .C(n6472), .Z(
        \CycleWaveform34[0] ) );
    GTECH_NAND2 U1500 ( .A(n6322), .B(n6472), .Z(n_168) );
    GTECH_AND2 U1501 ( .A(\*cell*469/U144/Z_0 ), .B(n6473), .Z(n_358) );
    GTECH_OAI21 U1502 ( .A(\IRQ[0] ), .B(n6474), .C(n6321), .Z(n_566) );
    GTECH_NAND2 U1503 ( .A(n6323), .B(n6321), .Z(n_565) );
    GTECH_NAND2 U1504 ( .A(n6475), .B(n6321), .Z(n_564) );
    GTECH_NOT U1505 ( .A(n6476), .Z(\IPRELOAD_Index3559[0] ) );
    GTECH_NAND2 U1506 ( .A(n6477), .B(n6478), .Z(\IPRELOAD_Index3559[1] ) );
    GTECH_NOT U1507 ( .A(n6479), .Z(\IPRELOAD_Index3559[2] ) );
    GTECH_NAND4 U1508 ( .A(n6480), .B(n6481), .C(n6482), .D(n6483), .Z(
        \IPRELOAD_Index3559[3] ) );
    GTECH_NAND2 U1509 ( .A(n6423), .B(n6322), .Z(\n2831[4][7][3] ) );
    GTECH_OAI21 U1510 ( .A(n6484), .B(n6471), .C(n6485), .Z(\n640[3] ) );
    GTECH_NOR3 U1511 ( .A(n6486), .B(n6487), .C(n6488), .Z(n6484) );
    GTECH_NAND3 U1512 ( .A(\NextInstruction[PARAMETER][3] ), .B(n6489), .C(
        \NextInstruction[PARAMETER][1] ), .Z(n6432) );
    GTECH_NAND3 U1513 ( .A(\NextInstruction[PARAMETER][0] ), .B(n6490), .C(
        \NextInstruction[PARAMETER][1] ), .Z(n6427) );
    GTECH_AOI222 U1514 ( .A(n6492), .B(n6322), .C(\Variables[0][-8][3]_wire ), 
        .D(n6493), .E(\sum2964[7] ), .F(n6494), .Z(n6491) );
    GTECH_AOI222 U1515 ( .A(n6496), .B(n6322), .C(\Variables[0][-8][2]_wire ), 
        .D(n6493), .E(\sum2964[6] ), .F(n6494), .Z(n6495) );
    GTECH_AOI222 U1516 ( .A(n6498), .B(n6322), .C(\Variables[0][-8][1]_wire ), 
        .D(n6493), .E(\sum2964[5] ), .F(n6494), .Z(n6497) );
    GTECH_AOI222 U1517 ( .A(n6500), .B(n6322), .C(\Variables[0][-8][0]_wire ), 
        .D(n6493), .E(\sum2964[4] ), .F(n6494), .Z(n6499) );
    GTECH_AOI222 U1518 ( .A(n6502), .B(n6322), .C(\Variables[0][-7][3]_wire ), 
        .D(n6493), .E(\sum2964[3] ), .F(n6494), .Z(n6501) );
    GTECH_AOI222 U1519 ( .A(n6504), .B(n6322), .C(\Variables[0][-7][2]_wire ), 
        .D(n6493), .E(\sum2964[2] ), .F(n6494), .Z(n6503) );
    GTECH_AOI222 U1520 ( .A(n6506), .B(n6322), .C(\Variables[0][-7][1]_wire ), 
        .D(n6493), .E(\sum2964[1] ), .F(n6494), .Z(n6505) );
    GTECH_AOI222 U1521 ( .A(n6508), .B(n6322), .C(\Variables[0][-7][0]_wire ), 
        .D(n6493), .E(\sum2964[0] ), .F(n6494), .Z(n6507) );
    GTECH_AOI222 U1522 ( .A(n6510), .B(n6322), .C(\Variables[0][-3][3]_wire ), 
        .D(n6511), .E(n6512), .F(\NextInstruction[PARAMETER][3] ), .Z(n6509)
         );
    GTECH_AOI222 U1523 ( .A(n6514), .B(n6322), .C(\Variables[0][-3][2]_wire ), 
        .D(n6511), .E(n6512), .F(\NextInstruction[PARAMETER][2] ), .Z(n6513)
         );
    GTECH_AOI222 U1524 ( .A(n6516), .B(n6322), .C(\Variables[0][-3][1]_wire ), 
        .D(n6511), .E(n6512), .F(\NextInstruction[PARAMETER][1] ), .Z(n6515)
         );
    GTECH_AOI222 U1525 ( .A(n6518), .B(n6322), .C(\Variables[0][-3][0]_wire ), 
        .D(n6511), .E(n6512), .F(\NextInstruction[PARAMETER][0] ), .Z(n6517)
         );
    GTECH_AND3 U1526 ( .A(n6520), .B(n6521), .C(n6522), .Z(n6519) );
    GTECH_AOI222 U1527 ( .A(n6523), .B(n6524), .C(n6525), .D(\sum2964[7] ), 
        .E(n6526), .F(\Variables[0][-8][3]_wire ), .Z(n6337) );
    GTECH_AOI222 U1528 ( .A(n6523), .B(n6527), .C(n6525), .D(\sum2964[6] ), 
        .E(n6526), .F(\Variables[0][-8][2]_wire ), .Z(n6338) );
    GTECH_AOI222 U1529 ( .A(n6523), .B(n6528), .C(n6525), .D(\sum2964[5] ), 
        .E(n6526), .F(\Variables[0][-8][1]_wire ), .Z(n6339) );
    GTECH_AOI222 U1530 ( .A(n6523), .B(n6529), .C(n6525), .D(\sum2964[4] ), 
        .E(n6526), .F(\Variables[0][-8][0]_wire ), .Z(n6340) );
    GTECH_AOI222 U1531 ( .A(n6523), .B(n6530), .C(n6525), .D(\sum2964[3] ), 
        .E(n6526), .F(\Variables[0][-7][3]_wire ), .Z(n6341) );
    GTECH_AOI222 U1532 ( .A(n6523), .B(n6531), .C(n6525), .D(\sum2964[2] ), 
        .E(n6526), .F(\Variables[0][-7][2]_wire ), .Z(n6342) );
    GTECH_AOI222 U1533 ( .A(n6523), .B(n6532), .C(n6525), .D(\sum2964[1] ), 
        .E(n6526), .F(\Variables[0][-7][1]_wire ), .Z(n6343) );
    GTECH_AOI222 U1534 ( .A(n6523), .B(n6533), .C(n6525), .D(\sum2964[0] ), 
        .E(n6526), .F(\Variables[0][-7][0]_wire ), .Z(n6344) );
    GTECH_AOI222 U1535 ( .A(n6523), .B(n6534), .C(n6535), .D(
        \NextInstruction[PARAMETER][3] ), .E(n6536), .F(
        \Variables[0][-3][3]_wire ), .Z(n6359) );
    GTECH_AOI222 U1536 ( .A(n6523), .B(n6537), .C(n6535), .D(
        \NextInstruction[PARAMETER][2] ), .E(n6536), .F(
        \Variables[0][-3][2]_wire ), .Z(n6360) );
    GTECH_AOI222 U1537 ( .A(n6523), .B(n6538), .C(n6535), .D(
        \NextInstruction[PARAMETER][1] ), .E(n6536), .F(
        \Variables[0][-3][1]_wire ), .Z(n6361) );
    GTECH_AOI222 U1538 ( .A(n6523), .B(n6539), .C(n6535), .D(
        \NextInstruction[PARAMETER][0] ), .E(n6536), .F(
        \Variables[0][-3][0]_wire ), .Z(n6362) );
    GTECH_AND8 U1539 ( .A(n6540), .B(n6541), .C(n6542), .D(n6543), .E(n6544), 
        .F(n6545), .G(n6546), .H(n6547), .Z(n6461) );
    GTECH_AND8 U1540 ( .A(n6548), .B(n6549), .C(n6550), .D(n6551), .E(n6552), 
        .F(n6553), .G(n6554), .H(n6555), .Z(n6464) );
    GTECH_AND8 U1541 ( .A(n6556), .B(n6557), .C(n6558), .D(n6559), .E(n6560), 
        .F(n6561), .G(n6562), .H(n6563), .Z(n6465) );
    GTECH_AND8 U1542 ( .A(n6564), .B(n6565), .C(n6566), .D(n6567), .E(n6568), 
        .F(n6569), .G(n6570), .H(n6571), .Z(n6466) );
    GTECH_AND8 U1543 ( .A(n6572), .B(n6573), .C(n6574), .D(n6575), .E(n6576), 
        .F(n6577), .G(n6578), .H(n6579), .Z(n6467) );
    GTECH_AND8 U1544 ( .A(n6580), .B(n6581), .C(n6582), .D(n6583), .E(n6584), 
        .F(n6585), .G(n6586), .H(n6587), .Z(n6468) );
    GTECH_AND8 U1545 ( .A(n6588), .B(n6589), .C(n6590), .D(n6591), .E(n6592), 
        .F(n6593), .G(n6594), .H(n6595), .Z(n6469) );
    GTECH_AND8 U1546 ( .A(n6596), .B(n6597), .C(n6598), .D(n6599), .E(n6600), 
        .F(n6601), .G(n6602), .H(n6603), .Z(n6470) );
    GTECH_AOI222 U1547 ( .A(\Interrupt_Index[2] ), .B(\IPRELOAD_Table3551[2] ), 
        .C(\Exception_Index[2] ), .D(n6604), .E(\IRQ_Index[2] ), .F(n6605), 
        .Z(n6479) );
    GTECH_AOI222 U1548 ( .A(\Interrupt_Index[0] ), .B(\IPRELOAD_Table3551[2] ), 
        .C(\Exception_Index[0] ), .D(n6604), .E(\IRQ_Index[0] ), .F(n6605), 
        .Z(n6476) );
    GTECH_OA21 U1549 ( .A(n6607), .B(n6608), .C(n6609), .Z(n6606) );
    GTECH_MAJ23 U1550 ( .A(n6611), .B(n6606), .C(n6612), .Z(n6610) );
    GTECH_OR2 U1551 ( .A(n6614), .B(n6615), .Z(n6613) );
    GTECH_AOI222 U1552 ( .A(n6431), .B(\Lower[3] ), .C(n6616), .D(n6617), .E(
        n6618), .F(n6619), .Z(n6433) );
    GTECH_AOI222 U1553 ( .A(n6431), .B(\Lower[2] ), .C(n6616), .D(n6620), .E(
        n6618), .F(n6621), .Z(n6436) );
    GTECH_AOI222 U1554 ( .A(n6431), .B(\Lower[1] ), .C(n6616), .D(n6622), .E(
        n6623), .F(n6618), .Z(n6437) );
    GTECH_AOI222 U1555 ( .A(n6431), .B(\Lower[0] ), .C(n6616), .D(n6624), .E(
        n6618), .F(n6625), .Z(n6438) );
    GTECH_OA21 U1556 ( .A(n6627), .B(n6628), .C(n6629), .Z(n6626) );
    GTECH_OA21 U1557 ( .A(n6628), .B(n6631), .C(n6632), .Z(n6630) );
    GTECH_AND3 U1558 ( .A(n6634), .B(n6450), .C(n6635), .Z(n6633) );
    GTECH_OR_NOT U1559 ( .A(MemoryReady), .B(n6636), .Z(n658) );
    GTECH_OAI2N2 U1560 ( .A(\Lower[3] ), .B(n6637), .C(n6491), .D(n6637), .Z(
        n6403) );
    GTECH_OAI2N2 U1561 ( .A(\Lower[2] ), .B(n6637), .C(n6495), .D(n6637), .Z(
        n6406) );
    GTECH_OAI2N2 U1562 ( .A(\Lower[1] ), .B(n6637), .C(n6497), .D(n6637), .Z(
        n6407) );
    GTECH_OAI2N2 U1563 ( .A(\Lower[0] ), .B(n6637), .C(n6499), .D(n6637), .Z(
        n6408) );
    GTECH_OAI2N2 U1564 ( .A(\Lower[3] ), .B(n6638), .C(n6501), .D(n6638), .Z(
        n6409) );
    GTECH_OAI2N2 U1565 ( .A(\Lower[2] ), .B(n6638), .C(n6503), .D(n6638), .Z(
        n6410) );
    GTECH_OAI2N2 U1566 ( .A(\Lower[1] ), .B(n6638), .C(n6505), .D(n6638), .Z(
        n6411) );
    GTECH_OAI2N2 U1567 ( .A(\Lower[0] ), .B(n6638), .C(n6507), .D(n6638), .Z(
        n6412) );
    GTECH_OAI2N2 U1568 ( .A(\Lower[3] ), .B(n6639), .C(n6509), .D(n6639), .Z(
        n6413) );
    GTECH_OAI2N2 U1569 ( .A(\Lower[2] ), .B(n6639), .C(n6513), .D(n6639), .Z(
        n6414) );
    GTECH_OAI2N2 U1570 ( .A(\Lower[1] ), .B(n6639), .C(n6515), .D(n6639), .Z(
        n6415) );
    GTECH_OAI2N2 U1571 ( .A(\Lower[0] ), .B(n6639), .C(n6517), .D(n6639), .Z(
        n6416) );
    GTECH_MUXI2 U1572 ( .A(n6641), .B(\IPRELOAD_Index[2] ), .S(n6642), .Z(
        n6640) );
    GTECH_XOR3 U1573 ( .A(n6335), .B(n6610), .C(n6643), .Z(n6619) );
    GTECH_XOR3 U1574 ( .A(n6612), .B(n6611), .C(n6644), .Z(n6621) );
    GTECH_OAI2N2 U1575 ( .A(n6645), .B(n6646), .C(n6645), .D(n6646), .Z(n6625)
         );
    GTECH_NOR3 U1576 ( .A(\IRQ[0] ), .B(\IRQ[2] ), .C(\IRQ[1] ), .Z(n6475) );
    GTECH_AND3 U1577 ( .A(n6647), .B(n6473), .C(IRQEnable), .Z(n_660) );
    GTECH_AND2 U1578 ( .A(n6648), .B(n6322), .Z(\IRQ2736[4] ) );
    GTECH_OR_NOT U1579 ( .A(n6649), .B(\IRQ[3] ), .Z(n6321) );
    GTECH_NAND3 U1580 ( .A(n6474), .B(n6325), .C(\IRQ[2] ), .Z(n6323) );
    GTECH_NOT U1581 ( .A(\IRQ[1] ), .Z(n6474) );
    GTECH_NOR3 U1582 ( .A(RegularJump), .B(ReturnJump), .C(InterruptJump), .Z(
        \IPRELOAD_Table3551[1] ) );
    GTECH_AND_NOT U1583 ( .A(\IPRELOAD_Table3551[1] ), .B(IRQJump), .Z(n6604)
         );
    GTECH_OA21 U1584 ( .A(IRQInProcess), .B(n7344), .C(n7341), .Z(n6328) );
    GTECH_AND_NOT U1585 ( .A(n6328), .B(\NextInstruction[INSTRUCTION][3] ), 
        .Z(n6650) );
    GTECH_NOT U1586 ( .A(\NextInstruction[INSTRUCTION][0] ), .Z(n6651) );
    GTECH_AND3 U1587 ( .A(n6650), .B(n6652), .C(
        \NextInstruction[INSTRUCTION][0] ), .Z(n6333) );
    GTECH_NOT U1588 ( .A(\NextInstruction[INSTRUCTION][2] ), .Z(n6627) );
    GTECH_AND3 U1589 ( .A(n6333), .B(n6628), .C(
        \NextInstruction[INSTRUCTION][2] ), .Z(\*cell*469/U12/Z_0 ) );
    GTECH_AND_NOT U1590 ( .A(n6336), .B(\NextInstruction[PARAMETER][2] ), .Z(
        n6490) );
    GTECH_NOT U1591 ( .A(\NextInstruction[PARAMETER][0] ), .Z(n6628) );
    GTECH_NOT U1592 ( .A(\NextInstruction[INSTRUCTION][1] ), .Z(n6652) );
    GTECH_AND3 U1593 ( .A(n6651), .B(n6627), .C(n6653), .Z(\*cell*469/U7/Z_0 )
         );
    GTECH_NOT U1594 ( .A(\NextInstruction[PARAMETER][3] ), .Z(n6336) );
    GTECH_NAND2 U1595 ( .A(\NextInstruction[PARAMETER][3] ), .B(n6655), .Z(
        n6654) );
    GTECH_NOT U1596 ( .A(\NextInstruction[INSTRUCTION][3] ), .Z(n6656) );
    GTECH_NAND4 U1597 ( .A(\NextInstruction[INSTRUCTION][3] ), .B(
        \NextInstruction[INSTRUCTION][0] ), .C(n6627), .D(n6652), .Z(n6657) );
    GTECH_AND_NOT U1598 ( .A(n6328), .B(n6657), .Z(n6329) );
    GTECH_AND_NOT U1599 ( .A(n6489), .B(n6654), .Z(n6460) );
    GTECH_NOT U1600 ( .A(\NextInstruction[PARAMETER][2] ), .Z(n6489) );
    GTECH_NAND3 U1601 ( .A(n6336), .B(n6655), .C(
        \NextInstruction[PARAMETER][2] ), .Z(n6658) );
    GTECH_NOT U1602 ( .A(\NextInstruction[PARAMETER][1] ), .Z(n6655) );
    GTECH_AND_NOT U1603 ( .A(\NextInstruction[PARAMETER][1] ), .B(n6489), .Z(
        n6659) );
    GTECH_AND_NOT U1604 ( .A(n6652), .B(\NextInstruction[INSTRUCTION][0] ), 
        .Z(n6660) );
    GTECH_NAND3 U1605 ( .A(n6651), .B(n6627), .C(
        \NextInstruction[INSTRUCTION][1] ), .Z(n6661) );
    GTECH_AND_NOT U1606 ( .A(n6656), .B(n6661), .Z(n6662) );
    GTECH_AND2 U1607 ( .A(n6490), .B(n6628), .Z(n6663) );
    GTECH_AND_NOT U1608 ( .A(n6322), .B(n6428), .Z(n6430) );
    GTECH_NAND2 U1609 ( .A(n6665), .B(n6666), .Z(n6664) );
    GTECH_AND_NOT U1610 ( .A(n6668), .B(n6664), .Z(n6667) );
    GTECH_NOR2 U1611 ( .A(n6656), .B(n6661), .Z(n6669) );
    GTECH_AND_NOT U1612 ( .A(n6670), .B(ResetStarted), .Z(n6435) );
    GTECH_NOR3 U1613 ( .A(ExceptionJump), .B(IRQJump), .C(ResetStarted), .Z(
        n6429) );
    GTECH_AND_NOT U1614 ( .A(n6462), .B(ResetStarted), .Z(n6463) );
    GTECH_NAND3 U1615 ( .A(n7347), .B(n7343), .C(n7342), .Z(n6671) );
    GTECH_AND_NOT U1616 ( .A(n6322), .B(n6671), .Z(n6424) );
    GTECH_AND_NOT U1617 ( .A(n6322), .B(OpCodeRegisterWrite), .Z(n6425) );
    GTECH_AND_NOT U1618 ( .A(n6663), .B(n6655), .Z(n6449) );
    GTECH_NOT U1619 ( .A(\gt_236/AEQB[2] ), .Z(n6520) );
    GTECH_NAND2 U1620 ( .A(n6322), .B(RegularRegisterWrite), .Z(n6672) );
    GTECH_NOR2 U1621 ( .A(n6673), .B(n6672), .Z(n6422) );
    GTECH_AND3 U1622 ( .A(n6522), .B(n6521), .C(\gt_236/AEQB[2] ), .Z(n6673)
         );
    GTECH_NAND2 U1623 ( .A(\RegularWriteRegister_Index[2] ), .B(
        \RegularWriteRegister_Index[1] ), .Z(n6674) );
    GTECH_OR_NOT U1624 ( .A(\RegularWriteRegister_Index[3] ), .B(
        \RegularWriteRegister_Index[0] ), .Z(n6675) );
    GTECH_NOT U1625 ( .A(\TableSelect[0] ), .Z(n6522) );
    GTECH_NOT U1626 ( .A(\TableSelect[1] ), .Z(n6521) );
    GTECH_AND3 U1627 ( .A(\TableSelect[0] ), .B(n6520), .C(\TableSelect[1] ), 
        .Z(n6676) );
    GTECH_AND3 U1628 ( .A(n6522), .B(n6520), .C(\TableSelect[1] ), .Z(n6677)
         );
    GTECH_AND3 U1629 ( .A(n6520), .B(n6521), .C(\TableSelect[0] ), .Z(n6678)
         );
    GTECH_NOR2 U1630 ( .A(n6680), .B(ResetStarted), .Z(n6679) );
    GTECH_NOT U1631 ( .A(\Lower[3] ), .Z(n6450) );
    GTECH_OR2 U1632 ( .A(n6675), .B(n6674), .Z(n6681) );
    GTECH_OR_NOT U1633 ( .A(n6423), .B(n6673), .Z(n6421) );
    GTECH_NOT U1634 ( .A(\Lower[2] ), .Z(n6453) );
    GTECH_NOT U1635 ( .A(\Lower[1] ), .Z(n6455) );
    GTECH_NOT U1636 ( .A(\Lower[0] ), .Z(n6456) );
    GTECH_OR2 U1637 ( .A(\RegularWriteRegister_Index[0] ), .B(
        \RegularWriteRegister_Index[3] ), .Z(n6682) );
    GTECH_AND_NOT U1638 ( .A(n6684), .B(ResetStarted), .Z(n6683) );
    GTECH_OR2 U1639 ( .A(n6682), .B(n6674), .Z(n6684) );
    GTECH_OR2 U1640 ( .A(\RegularWriteRegister_Index[1] ), .B(n6686), .Z(n6685
        ) );
    GTECH_NOR2 U1641 ( .A(ResetStarted), .B(n6688), .Z(n6687) );
    GTECH_NOR2 U1642 ( .A(n6675), .B(n6685), .Z(n6688) );
    GTECH_NOR2 U1643 ( .A(ResetStarted), .B(n6690), .Z(n6689) );
    GTECH_NOR2 U1644 ( .A(n6682), .B(n6685), .Z(n6690) );
    GTECH_NAND2 U1645 ( .A(n6686), .B(\RegularWriteRegister_Index[1] ), .Z(
        n6691) );
    GTECH_AND2 U1646 ( .A(n6693), .B(n6322), .Z(n6692) );
    GTECH_OR2 U1647 ( .A(n6691), .B(n6675), .Z(n6693) );
    GTECH_AND_NOT U1648 ( .A(n6695), .B(ResetStarted), .Z(n6694) );
    GTECH_OR2 U1649 ( .A(n6691), .B(n6682), .Z(n6695) );
    GTECH_NOR2 U1650 ( .A(\RegularWriteRegister_Index[2] ), .B(
        \RegularWriteRegister_Index[1] ), .Z(n6696) );
    GTECH_NOR2 U1651 ( .A(ResetStarted), .B(n6698), .Z(n6697) );
    GTECH_AND_NOT U1652 ( .A(n6696), .B(n6675), .Z(n6698) );
    GTECH_NOR2 U1653 ( .A(ResetStarted), .B(n6700), .Z(n6699) );
    GTECH_AND_NOT U1654 ( .A(n6696), .B(n6682), .Z(n6700) );
    GTECH_OR_NOT U1655 ( .A(\RegularWriteRegister_Index[0] ), .B(
        \RegularWriteRegister_Index[3] ), .Z(n6701) );
    GTECH_AND2 U1656 ( .A(n6424), .B(n6519), .Z(n6493) );
    GTECH_AND2 U1657 ( .A(n6671), .B(n6519), .Z(n6494) );
    GTECH_AND2 U1658 ( .A(\RegularWriteRegister_Index[0] ), .B(
        \RegularWriteRegister_Index[3] ), .Z(n6702) );
    GTECH_AND2 U1659 ( .A(n6704), .B(n6322), .Z(n6703) );
    GTECH_OR2 U1660 ( .A(n6701), .B(n6691), .Z(n6704) );
    GTECH_NOR2 U1661 ( .A(ResetStarted), .B(n6706), .Z(n6705) );
    GTECH_AND_NOT U1662 ( .A(n6702), .B(n6691), .Z(n6706) );
    GTECH_AND2 U1663 ( .A(n6708), .B(n6322), .Z(n6707) );
    GTECH_OR2 U1664 ( .A(n6701), .B(n6685), .Z(n6708) );
    GTECH_AND2 U1665 ( .A(n6425), .B(n6519), .Z(n6511) );
    GTECH_AND2 U1666 ( .A(OpCodeRegisterWrite), .B(n6519), .Z(n6512) );
    GTECH_NOR2 U1667 ( .A(ResetStarted), .B(n6710), .Z(n6709) );
    GTECH_NOR2 U1668 ( .A(n6701), .B(n6674), .Z(n6710) );
    GTECH_OR_NOT U1669 ( .A(n6712), .B(n6322), .Z(n6711) );
    GTECH_AND_NOT U1670 ( .A(n6702), .B(n6674), .Z(n6712) );
    GTECH_NOR2 U1671 ( .A(n6672), .B(n6676), .Z(n6420) );
    GTECH_OR_NOT U1672 ( .A(n6423), .B(n6676), .Z(n6419) );
    GTECH_NOR2 U1673 ( .A(n6677), .B(n6672), .Z(n6418) );
    GTECH_OR_NOT U1674 ( .A(n6423), .B(n6677), .Z(n6417) );
    GTECH_NOR2 U1675 ( .A(n6678), .B(n6672), .Z(n6405) );
    GTECH_OR_NOT U1676 ( .A(n6423), .B(n6678), .Z(n6404) );
    GTECH_NOR2 U1677 ( .A(n6519), .B(n6672), .Z(n6347) );
    GTECH_NOR2 U1678 ( .A(n6713), .B(n6423), .Z(n6523) );
    GTECH_OA21 U1679 ( .A(n6713), .B(n6423), .C(n6671), .Z(n6525) );
    GTECH_AND3 U1680 ( .A(n6424), .B(n6713), .C(RegularRegisterWrite), .Z(
        n6526) );
    GTECH_OA21 U1681 ( .A(n6713), .B(n6423), .C(OpCodeRegisterWrite), .Z(n6535
        ) );
    GTECH_AND3 U1682 ( .A(n6425), .B(n6713), .C(RegularRegisterWrite), .Z(
        n6536) );
    GTECH_NAND2 U1683 ( .A(n6322), .B(\NextInstruction[INSTRUCTION][1] ), .Z(
        n6451) );
    GTECH_NOT U1684 ( .A(\Upper[3] ), .Z(n6714) );
    GTECH_NOT U1685 ( .A(\Upper[2] ), .Z(n6715) );
    GTECH_NOT U1686 ( .A(\Upper[1] ), .Z(n6716) );
    GTECH_AND3 U1687 ( .A(n6490), .B(n6655), .C(
        \NextInstruction[PARAMETER][0] ), .Z(n6448) );
    GTECH_NOT U1688 ( .A(\IPRELOAD_Index[2] ), .Z(n6641) );
    GTECH_NOT U1689 ( .A(\add_417/carry[1] ), .Z(n6717) );
    GTECH_AND_NOT U1690 ( .A(\IPRELOAD_Index[1] ), .B(n6717), .Z(n6642) );
    GTECH_AND2 U1691 ( .A(n6719), .B(\IPRELOAD_Index[2] ), .Z(n6718) );
    GTECH_NOT U1692 ( .A(\IPRELOAD_Table[2] ), .Z(n6720) );
    GTECH_AND3 U1693 ( .A(n6722), .B(n6723), .C(\IPRELOAD_Table[2] ), .Z(n6721
        ) );
    GTECH_NOT U1694 ( .A(\IPRELOAD_Table[0] ), .Z(n6722) );
    GTECH_NOT U1695 ( .A(\IPRELOAD_Table[1] ), .Z(n6723) );
    GTECH_AND3 U1696 ( .A(\IPRELOAD_Table[0] ), .B(n6720), .C(
        \IPRELOAD_Table[1] ), .Z(n6724) );
    GTECH_AND3 U1697 ( .A(n6722), .B(n6720), .C(\IPRELOAD_Table[1] ), .Z(n6725
        ) );
    GTECH_NOR3 U1698 ( .A(\IPRELOAD_Table[1] ), .B(\IPRELOAD_Table[2] ), .C(
        n6722), .Z(n6726) );
    GTECH_AND3 U1699 ( .A(n6723), .B(n6720), .C(n6722), .Z(n6727) );
    GTECH_NAND2 U1700 ( .A(n6718), .B(n6642), .Z(n6728) );
    GTECH_AND_NOT U1701 ( .A(\IPRELOAD_Index[1] ), .B(\add_417/carry[1] ), .Z(
        n6729) );
    GTECH_NAND2 U1702 ( .A(n6718), .B(n6729), .Z(n6730) );
    GTECH_OR2 U1703 ( .A(\IPRELOAD_Index[1] ), .B(n6717), .Z(n6731) );
    GTECH_OR_NOT U1704 ( .A(n6731), .B(n6718), .Z(n6732) );
    GTECH_OR2 U1705 ( .A(\IPRELOAD_Index[1] ), .B(\add_417/carry[1] ), .Z(
        n6733) );
    GTECH_AND_NOT U1706 ( .A(n6718), .B(n6733), .Z(n6734) );
    GTECH_OR_NOT U1707 ( .A(\IPRELOAD_Index[2] ), .B(n6719), .Z(n6735) );
    GTECH_OR_NOT U1708 ( .A(n6735), .B(n6642), .Z(n6736) );
    GTECH_AND_NOT U1709 ( .A(n6729), .B(n6735), .Z(n6737) );
    GTECH_OR2 U1710 ( .A(n6735), .B(n6731), .Z(n6738) );
    GTECH_NOR2 U1711 ( .A(n6735), .B(n6733), .Z(n6739) );
    GTECH_NOT U1712 ( .A(\IPRELOAD_Index[3] ), .Z(n6719) );
    GTECH_OR_NOT U1713 ( .A(n6641), .B(\IPRELOAD_Index[3] ), .Z(n6740) );
    GTECH_OR_NOT U1714 ( .A(n6740), .B(n6642), .Z(n6741) );
    GTECH_AND_NOT U1715 ( .A(n6729), .B(n6740), .Z(n6742) );
    GTECH_OR2 U1716 ( .A(n6740), .B(n6731), .Z(n6743) );
    GTECH_NOR2 U1717 ( .A(n6733), .B(n6740), .Z(n6744) );
    GTECH_OR_NOT U1718 ( .A(n6719), .B(n6641), .Z(n6745) );
    GTECH_OR_NOT U1719 ( .A(n6745), .B(n6642), .Z(n6746) );
    GTECH_OR_NOT U1720 ( .A(n6745), .B(n6729), .Z(n6747) );
    GTECH_OR2 U1721 ( .A(n6731), .B(n6745), .Z(n6748) );
    GTECH_OR2 U1722 ( .A(n6733), .B(n6745), .Z(n6749) );
    GTECH_NOT U1723 ( .A(Condition), .Z(n6462) );
    GTECH_OA21 U1724 ( .A(n6642), .B(n6719), .C(n6751), .Z(n6750) );
    GTECH_OR_NOT U1725 ( .A(n6753), .B(n6750), .Z(n6752) );
    GTECH_NAND2 U1726 ( .A(n6717), .B(n6640), .Z(n6754) );
    GTECH_OR2 U1727 ( .A(n6752), .B(n6754), .Z(n6755) );
    GTECH_OR_NOT U1728 ( .A(n6717), .B(n6640), .Z(n6756) );
    GTECH_OR2 U1729 ( .A(n6756), .B(n6752), .Z(n6757) );
    GTECH_AND_NOT U1730 ( .A(n6731), .B(n6729), .Z(n6753) );
    GTECH_AND_NOT U1731 ( .A(n6750), .B(n6759), .Z(n6758) );
    GTECH_OR_NOT U1732 ( .A(n6754), .B(n6758), .Z(n6760) );
    GTECH_AND_NOT U1733 ( .A(n6758), .B(n6756), .Z(n6761) );
    GTECH_OR_NOT U1734 ( .A(n6640), .B(n6717), .Z(n6762) );
    GTECH_OR2 U1735 ( .A(n6752), .B(n6762), .Z(n6763) );
    GTECH_OR_NOT U1736 ( .A(n6640), .B(\add_417/carry[1] ), .Z(n6764) );
    GTECH_NOR2 U1737 ( .A(n6752), .B(n6764), .Z(n6765) );
    GTECH_OR_NOT U1738 ( .A(n6762), .B(n6758), .Z(n6766) );
    GTECH_AND_NOT U1739 ( .A(n6758), .B(n6764), .Z(n6767) );
    GTECH_OR2 U1740 ( .A(n6750), .B(n6753), .Z(n6768) );
    GTECH_OR2 U1741 ( .A(n6768), .B(n6754), .Z(n6769) );
    GTECH_NOR2 U1742 ( .A(n6756), .B(n6768), .Z(n6770) );
    GTECH_OR2 U1743 ( .A(n6750), .B(n6759), .Z(n6771) );
    GTECH_OR2 U1744 ( .A(n6771), .B(n6754), .Z(n6772) );
    GTECH_NOR2 U1745 ( .A(n6756), .B(n6771), .Z(n6773) );
    GTECH_OR2 U1746 ( .A(n6762), .B(n6768), .Z(n6774) );
    GTECH_NOR2 U1747 ( .A(n6764), .B(n6768), .Z(n6775) );
    GTECH_OR2 U1748 ( .A(n6762), .B(n6771), .Z(n6776) );
    GTECH_OR2 U1749 ( .A(n6764), .B(n6771), .Z(n6777) );
    GTECH_AND_NOT U1750 ( .A(n6628), .B(n6432), .Z(n6431) );
    GTECH_AND2 U1751 ( .A(IRQJump), .B(\IPRELOAD_Table3551[1] ), .Z(n6605) );
    GTECH_AND3 U1752 ( .A(n6480), .B(n6481), .C(InterruptJump), .Z(
        \IPRELOAD_Table3551[2] ) );
    GTECH_NOT U1753 ( .A(RegularJump), .Z(n6480) );
    GTECH_OR_NOT U1754 ( .A(ResetStarted), .B(n6471), .Z(n6426) );
    GTECH_NOT U1755 ( .A(MemoryReadValue[3]), .Z(n6440) );
    GTECH_AND2 U1756 ( .A(n6449), .B(n6662), .Z(n6778) );
    GTECH_AND_NOT U1757 ( .A(n6663), .B(\NextInstruction[PARAMETER][1] ), .Z(
        n6635) );
    GTECH_AND2 U1758 ( .A(\Upper[0] ), .B(\Upper[2] ), .Z(n6779) );
    GTECH_NAND2 U1759 ( .A(\Upper[3] ), .B(n6716), .Z(n6780) );
    GTECH_NAND2 U1760 ( .A(n6781), .B(n6782), .Z(n6510) );
    GTECH_OR_NOT U1761 ( .A(n6780), .B(n6779), .Z(n6783) );
    GTECH_NOR2 U1762 ( .A(n6785), .B(\Upper[2] ), .Z(n6784) );
    GTECH_NAND2 U1763 ( .A(n6786), .B(n6787), .Z(n6502) );
    GTECH_NOR2 U1764 ( .A(n6789), .B(n6780), .Z(n6788) );
    GTECH_AND_NOT U1765 ( .A(n6785), .B(\Upper[2] ), .Z(n6790) );
    GTECH_NAND2 U1766 ( .A(n6791), .B(n6792), .Z(n6492) );
    GTECH_OR_NOT U1767 ( .A(n6780), .B(n6790), .Z(n6793) );
    GTECH_NAND2 U1768 ( .A(\Upper[1] ), .B(n6714), .Z(n6794) );
    GTECH_AND_NOT U1769 ( .A(n6779), .B(n6794), .Z(n6795) );
    GTECH_AND_NOT U1770 ( .A(n6785), .B(n6715), .Z(n6796) );
    GTECH_AND_NOT U1771 ( .A(n6796), .B(n6794), .Z(n6797) );
    GTECH_NAND2 U1772 ( .A(n6714), .B(n6716), .Z(n6798) );
    GTECH_AND_NOT U1773 ( .A(n6779), .B(n6798), .Z(n6799) );
    GTECH_AND_NOT U1774 ( .A(n6796), .B(n6798), .Z(n6800) );
    GTECH_AND_NOT U1775 ( .A(n6784), .B(n6794), .Z(n6801) );
    GTECH_AND_NOT U1776 ( .A(n6790), .B(n6794), .Z(n6802) );
    GTECH_AND_NOT U1777 ( .A(n6784), .B(n6798), .Z(n6803) );
    GTECH_AND_NOT U1778 ( .A(n6790), .B(n6798), .Z(n6804) );
    GTECH_NAND2 U1779 ( .A(\Upper[1] ), .B(\Upper[3] ), .Z(n6805) );
    GTECH_OR_NOT U1780 ( .A(n6805), .B(n6779), .Z(n6806) );
    GTECH_AND_NOT U1781 ( .A(n6796), .B(n6805), .Z(n6807) );
    GTECH_AND_NOT U1782 ( .A(n6796), .B(n6780), .Z(n6808) );
    GTECH_NOR2 U1783 ( .A(n6789), .B(n6805), .Z(n6809) );
    GTECH_AND_NOT U1784 ( .A(n6790), .B(n6805), .Z(n6810) );
    GTECH_AND2 U1785 ( .A(n6635), .B(n6662), .Z(n6811) );
    GTECH_OR_NOT U1786 ( .A(\NextInstruction[PARAMETER][3] ), .B(\Lower[3] ), 
        .Z(n6631) );
    GTECH_AND_NOT U1787 ( .A(\NextInstruction[PARAMETER][0] ), .B(n6658), .Z(
        n6812) );
    GTECH_AND_NOT U1788 ( .A(n6813), .B(n6814), .Z(n6607) );
    GTECH_NAND2 U1789 ( .A(\Upper[1] ), .B(n6336), .Z(n6815) );
    GTECH_OR_NOT U1790 ( .A(n6646), .B(n6645), .Z(n6608) );
    GTECH_OAI21 U1791 ( .A(n6607), .B(n6608), .C(n6609), .Z(n6644) );
    GTECH_AND_NOT U1792 ( .A(n6816), .B(n6817), .Z(n6611) );
    GTECH_NAND2 U1793 ( .A(n6336), .B(\Upper[2] ), .Z(n6612) );
    GTECH_NOR2 U1794 ( .A(n6628), .B(n6432), .Z(n6818) );
    GTECH_NOR2 U1795 ( .A(\NextInstruction[PARAMETER][0] ), .B(n6658), .Z(
        n6332) );
    GTECH_AND4 U1796 ( .A(\NextInstruction[INSTRUCTION][1] ), .B(
        \NextInstruction[INSTRUCTION][2] ), .C(n6651), .D(n6656), .Z(n6486) );
    GTECH_OR3 U1797 ( .A(n6654), .B(n6628), .C(n6489), .Z(n6819) );
    GTECH_AND2 U1798 ( .A(n6460), .B(\NextInstruction[PARAMETER][0] ), .Z(
        n6820) );
    GTECH_NAND2 U1799 ( .A(n6628), .B(n6460), .Z(n6821) );
    GTECH_NOR3 U1800 ( .A(n6628), .B(\NextInstruction[PARAMETER][3] ), .C(
        n6665), .Z(n6330) );
    GTECH_AND3 U1801 ( .A(n6336), .B(n6628), .C(n6659), .Z(n6822) );
    GTECH_OR3 U1802 ( .A(n6336), .B(n6628), .C(n6665), .Z(n6823) );
    GTECH_NOR3 U1803 ( .A(n6336), .B(\NextInstruction[PARAMETER][0] ), .C(
        n6665), .Z(n6824) );
    GTECH_NOR3 U1804 ( .A(n6654), .B(\NextInstruction[PARAMETER][0] ), .C(
        n6489), .Z(n6618) );
    GTECH_AND3 U1805 ( .A(\NextInstruction[INSTRUCTION][3] ), .B(n6627), .C(
        n6660), .Z(n6487) );
    GTECH_NAND2 U1806 ( .A(n6322), .B(n6328), .Z(n6825) );
    GTECH_NOT U1807 ( .A(MemoryReadValue[2]), .Z(n6442) );
    GTECH_NAND2 U1808 ( .A(n6826), .B(n6827), .Z(n6514) );
    GTECH_NAND2 U1809 ( .A(n6828), .B(n6829), .Z(n6504) );
    GTECH_NAND2 U1810 ( .A(n6830), .B(n6831), .Z(n6496) );
    GTECH_NAND2 U1811 ( .A(n6336), .B(\Lower[2] ), .Z(n6816) );
    GTECH_NOT U1812 ( .A(MemoryReadValue[1]), .Z(n6444) );
    GTECH_NAND2 U1813 ( .A(n6832), .B(n6833), .Z(n6516) );
    GTECH_NAND2 U1814 ( .A(n6834), .B(n6835), .Z(n6506) );
    GTECH_NAND2 U1815 ( .A(n6836), .B(n6837), .Z(n6498) );
    GTECH_NAND2 U1816 ( .A(\Lower[1] ), .B(n6336), .Z(n6813) );
    GTECH_NOT U1817 ( .A(MemoryReadValue[0]), .Z(n6446) );
    GTECH_NAND2 U1818 ( .A(n6838), .B(n6839), .Z(n6518) );
    GTECH_NAND2 U1819 ( .A(n6840), .B(n6841), .Z(n6508) );
    GTECH_NAND2 U1820 ( .A(n6842), .B(n6843), .Z(n6500) );
    GTECH_OR2 U1821 ( .A(n6825), .B(n6844), .Z(n6434) );
    GTECH_AND_NOT U1822 ( .A(n6336), .B(\Lower[0] ), .Z(n6615) );
    GTECH_AND_NOT U1823 ( .A(n6845), .B(n6657), .Z(n6331) );
    GTECH_MUX2 U1824 ( .A(\NextInstruction[PARAMETER][3] ), .B(\Upper[3] ), 
        .S(\NextInstruction[INSTRUCTION][1] ), .Z(
        \RegularWriteRegister_Index848[3] ) );
    GTECH_MUX2 U1825 ( .A(\NextInstruction[PARAMETER][2] ), .B(\Upper[2] ), 
        .S(\NextInstruction[INSTRUCTION][1] ), .Z(
        \RegularWriteRegister_Index848[2] ) );
    GTECH_MUX2 U1826 ( .A(\NextInstruction[PARAMETER][1] ), .B(\Upper[1] ), 
        .S(\NextInstruction[INSTRUCTION][1] ), .Z(
        \RegularWriteRegister_Index848[1] ) );
    GTECH_MUX2 U1827 ( .A(\NextInstruction[PARAMETER][0] ), .B(\Upper[0] ), 
        .S(\NextInstruction[INSTRUCTION][1] ), .Z(
        \RegularWriteRegister_Index848[0] ) );
    GTECH_MUX2 U1828 ( .A(\Variables[0][-2][3]_wire ), .B(\Upper[3] ), .S(
        Write_wire), .Z(\MemoryPtr3672[7] ) );
    GTECH_MUX2 U1829 ( .A(\Variables[0][-2][2]_wire ), .B(\Upper[2] ), .S(
        Write_wire), .Z(\MemoryPtr3672[6] ) );
    GTECH_MUX2 U1830 ( .A(\Variables[0][-2][1]_wire ), .B(\Upper[1] ), .S(
        Write_wire), .Z(\MemoryPtr3672[5] ) );
    GTECH_MUX2 U1831 ( .A(\Variables[0][-2][0]_wire ), .B(\Upper[0] ), .S(
        Write_wire), .Z(\MemoryPtr3672[4] ) );
    GTECH_MUX2 U1832 ( .A(\Variables[0][-1][3]_wire ), .B(\Lower[3] ), .S(
        Write_wire), .Z(\MemoryPtr3672[3] ) );
    GTECH_MUX2 U1833 ( .A(\Variables[0][-1][2]_wire ), .B(\Lower[2] ), .S(
        Write_wire), .Z(\MemoryPtr3672[2] ) );
    GTECH_MUX2 U1834 ( .A(\Lower[1] ), .B(\Variables[0][-1][1]_wire ), .S(
        n6317), .Z(\MemoryPtr3672[1] ) );
    GTECH_MUX2 U1835 ( .A(\Lower[0] ), .B(\Variables[0][-1][0]_wire ), .S(
        n6317), .Z(\MemoryPtr3672[0] ) );
    GTECH_AOI2N2 U1836 ( .A(n6846), .B(n6627), .C(
        \NextInstruction[INSTRUCTION][3] ), .D(n6627), .Z(n6326) );
    GTECH_AND5 U1837 ( .A(net109), .B(net112), .C(net108), .D(net111), .E(
        net110), .Z(n6847) );
    GTECH_OA21 U1838 ( .A(n6448), .B(n6652), .C(n6650), .Z(n6653) );
    GTECH_OA21 U1839 ( .A(\NextInstruction[PARAMETER][0] ), .B(n6336), .C(
        n6654), .Z(n6668) );
    GTECH_AO22 U1840 ( .A(n6662), .B(n6663), .C(n6667), .D(n6669), .Z(n6488)
         );
    GTECH_AOI21 U1841 ( .A(MemoryReady), .B(Read_wire), .C(ResetStarted), .Z(
        n6485) );
    GTECH_AOI222 U1842 ( .A(n6677), .B(\Variables[2][7][3]_wire ), .C(n6673), 
        .D(\Variables[4][7][3]_wire ), .E(n6676), .F(\Variables[3][7][3]_wire 
        ), .Z(n6848) );
    GTECH_AOI22 U1843 ( .A(n6519), .B(\Variables[0][7][3]_wire ), .C(
        \Variables[1][7][3]_wire ), .D(n6678), .Z(n6849) );
    GTECH_AOI222 U1844 ( .A(\Variables[2][7][2]_wire ), .B(n6677), .C(
        \Variables[4][7][2]_wire ), .D(n6673), .E(\Variables[3][7][2]_wire ), 
        .F(n6676), .Z(n6850) );
    GTECH_AOI22 U1845 ( .A(n6519), .B(\Variables[0][7][2]_wire ), .C(n6678), 
        .D(\Variables[1][7][2]_wire ), .Z(n6851) );
    GTECH_AOI222 U1846 ( .A(\Variables[2][7][1]_wire ), .B(n6677), .C(
        \Variables[4][7][1]_wire ), .D(n6673), .E(\Variables[3][7][1]_wire ), 
        .F(n6676), .Z(n6852) );
    GTECH_AOI22 U1847 ( .A(n6519), .B(\Variables[0][7][1]_wire ), .C(n6678), 
        .D(\Variables[1][7][1]_wire ), .Z(n6853) );
    GTECH_AOI222 U1848 ( .A(\Variables[2][7][0]_wire ), .B(n6677), .C(
        \Variables[4][7][0]_wire ), .D(n6673), .E(\Variables[3][7][0]_wire ), 
        .F(n6676), .Z(n6854) );
    GTECH_AOI22 U1849 ( .A(n6519), .B(\Variables[0][7][0]_wire ), .C(n6678), 
        .D(\Variables[1][7][0]_wire ), .Z(n6855) );
    GTECH_AOI222 U1850 ( .A(\Variables[2][6][3]_wire ), .B(n6677), .C(
        \Variables[4][6][3]_wire ), .D(n6673), .E(\Variables[3][6][3]_wire ), 
        .F(n6676), .Z(n6856) );
    GTECH_AOI22 U1851 ( .A(n6519), .B(\Variables[0][6][3]_wire ), .C(n6678), 
        .D(\Variables[1][6][3]_wire ), .Z(n6857) );
    GTECH_AOI222 U1852 ( .A(\Variables[2][6][2]_wire ), .B(n6677), .C(
        \Variables[4][6][2]_wire ), .D(n6673), .E(\Variables[3][6][2]_wire ), 
        .F(n6676), .Z(n6858) );
    GTECH_AOI22 U1853 ( .A(n6519), .B(\Variables[0][6][2]_wire ), .C(n6678), 
        .D(\Variables[1][6][2]_wire ), .Z(n6859) );
    GTECH_AOI222 U1854 ( .A(\Variables[2][6][1]_wire ), .B(n6677), .C(
        \Variables[4][6][1]_wire ), .D(n6673), .E(\Variables[3][6][1]_wire ), 
        .F(n6676), .Z(n6860) );
    GTECH_AOI22 U1855 ( .A(n6519), .B(\Variables[0][6][1]_wire ), .C(n6678), 
        .D(\Variables[1][6][1]_wire ), .Z(n6861) );
    GTECH_AOI222 U1856 ( .A(\Variables[2][6][0]_wire ), .B(n6677), .C(
        \Variables[4][6][0]_wire ), .D(n6673), .E(\Variables[3][6][0]_wire ), 
        .F(n6676), .Z(n6862) );
    GTECH_AOI22 U1857 ( .A(n6678), .B(\Variables[1][6][0]_wire ), .C(n6519), 
        .D(\Variables[0][6][0]_wire ), .Z(n6863) );
    GTECH_AOI222 U1858 ( .A(\Variables[2][5][3]_wire ), .B(n6677), .C(
        \Variables[4][5][3]_wire ), .D(n6673), .E(\Variables[3][5][3]_wire ), 
        .F(n6676), .Z(n6864) );
    GTECH_AOI22 U1859 ( .A(n6519), .B(\Variables[0][5][3]_wire ), .C(n6678), 
        .D(\Variables[1][5][3]_wire ), .Z(n6865) );
    GTECH_AOI222 U1860 ( .A(\Variables[2][5][2]_wire ), .B(n6677), .C(
        \Variables[4][5][2]_wire ), .D(n6673), .E(\Variables[3][5][2]_wire ), 
        .F(n6676), .Z(n6866) );
    GTECH_AOI22 U1861 ( .A(n6519), .B(\Variables[0][5][2]_wire ), .C(n6678), 
        .D(\Variables[1][5][2]_wire ), .Z(n6867) );
    GTECH_AOI222 U1862 ( .A(\Variables[2][5][1]_wire ), .B(n6677), .C(
        \Variables[4][5][1]_wire ), .D(n6673), .E(\Variables[3][5][1]_wire ), 
        .F(n6676), .Z(n6868) );
    GTECH_AOI22 U1863 ( .A(n6519), .B(\Variables[0][5][1]_wire ), .C(n6678), 
        .D(\Variables[1][5][1]_wire ), .Z(n6869) );
    GTECH_AOI222 U1864 ( .A(\Variables[2][5][0]_wire ), .B(n6677), .C(
        \Variables[4][5][0]_wire ), .D(n6673), .E(\Variables[3][5][0]_wire ), 
        .F(n6676), .Z(n6870) );
    GTECH_AOI22 U1865 ( .A(n6519), .B(\Variables[0][5][0]_wire ), .C(n6678), 
        .D(\Variables[1][5][0]_wire ), .Z(n6871) );
    GTECH_AOI222 U1866 ( .A(\Variables[2][4][3]_wire ), .B(n6677), .C(
        \Variables[4][4][3]_wire ), .D(n6673), .E(\Variables[3][4][3]_wire ), 
        .F(n6676), .Z(n6872) );
    GTECH_AOI22 U1867 ( .A(n6519), .B(\Variables[0][4][3]_wire ), .C(n6678), 
        .D(\Variables[1][4][3]_wire ), .Z(n6873) );
    GTECH_AOI222 U1868 ( .A(\Variables[2][4][2]_wire ), .B(n6677), .C(
        \Variables[4][4][2]_wire ), .D(n6673), .E(\Variables[3][4][2]_wire ), 
        .F(n6676), .Z(n6874) );
    GTECH_AOI22 U1869 ( .A(n6519), .B(\Variables[0][4][2]_wire ), .C(n6678), 
        .D(\Variables[1][4][2]_wire ), .Z(n6875) );
    GTECH_AOI222 U1870 ( .A(\Variables[2][4][1]_wire ), .B(n6677), .C(
        \Variables[4][4][1]_wire ), .D(n6673), .E(\Variables[3][4][1]_wire ), 
        .F(n6676), .Z(n6876) );
    GTECH_AOI22 U1871 ( .A(n6519), .B(\Variables[0][4][1]_wire ), .C(n6678), 
        .D(\Variables[1][4][1]_wire ), .Z(n6877) );
    GTECH_AOI222 U1872 ( .A(\Variables[2][4][0]_wire ), .B(n6677), .C(
        \Variables[4][4][0]_wire ), .D(n6673), .E(\Variables[3][4][0]_wire ), 
        .F(n6676), .Z(n6878) );
    GTECH_AOI22 U1873 ( .A(n6519), .B(\Variables[0][4][0]_wire ), .C(n6678), 
        .D(\Variables[1][4][0]_wire ), .Z(n6879) );
    GTECH_AOI222 U1874 ( .A(\Variables[2][3][3]_wire ), .B(n6677), .C(
        \Variables[4][3][3]_wire ), .D(n6673), .E(\Variables[3][3][3]_wire ), 
        .F(n6676), .Z(n6880) );
    GTECH_AOI22 U1875 ( .A(n6519), .B(\Variables[0][3][3]_wire ), .C(n6678), 
        .D(\Variables[1][3][3]_wire ), .Z(n6881) );
    GTECH_AOI222 U1876 ( .A(\Variables[2][3][2]_wire ), .B(n6677), .C(
        \Variables[4][3][2]_wire ), .D(n6673), .E(\Variables[3][3][2]_wire ), 
        .F(n6676), .Z(n6882) );
    GTECH_AOI22 U1877 ( .A(n6519), .B(\Variables[0][3][2]_wire ), .C(n6678), 
        .D(\Variables[1][3][2]_wire ), .Z(n6883) );
    GTECH_AOI222 U1878 ( .A(\Variables[2][3][1]_wire ), .B(n6677), .C(
        \Variables[4][3][1]_wire ), .D(n6673), .E(\Variables[3][3][1]_wire ), 
        .F(n6676), .Z(n6884) );
    GTECH_AOI22 U1879 ( .A(n6519), .B(\Variables[0][3][1]_wire ), .C(n6678), 
        .D(\Variables[1][3][1]_wire ), .Z(n6885) );
    GTECH_AOI222 U1880 ( .A(\Variables[2][3][0]_wire ), .B(n6677), .C(
        \Variables[4][3][0]_wire ), .D(n6673), .E(\Variables[3][3][0]_wire ), 
        .F(n6676), .Z(n6886) );
    GTECH_AOI22 U1881 ( .A(n6519), .B(\Variables[0][3][0]_wire ), .C(n6678), 
        .D(\Variables[1][3][0]_wire ), .Z(n6887) );
    GTECH_AOI222 U1882 ( .A(\Variables[2][2][3]_wire ), .B(n6677), .C(
        \Variables[4][2][3]_wire ), .D(n6673), .E(\Variables[3][2][3]_wire ), 
        .F(n6676), .Z(n6888) );
    GTECH_AOI22 U1883 ( .A(n6519), .B(\Variables[0][2][3]_wire ), .C(n6678), 
        .D(\Variables[1][2][3]_wire ), .Z(n6889) );
    GTECH_AOI222 U1884 ( .A(\Variables[2][2][2]_wire ), .B(n6677), .C(
        \Variables[4][2][2]_wire ), .D(n6673), .E(\Variables[3][2][2]_wire ), 
        .F(n6676), .Z(n6890) );
    GTECH_AOI22 U1885 ( .A(n6519), .B(\Variables[0][2][2]_wire ), .C(n6678), 
        .D(\Variables[1][2][2]_wire ), .Z(n6891) );
    GTECH_AOI222 U1886 ( .A(\Variables[2][2][1]_wire ), .B(n6677), .C(
        \Variables[4][2][1]_wire ), .D(n6673), .E(\Variables[3][2][1]_wire ), 
        .F(n6676), .Z(n6892) );
    GTECH_AOI22 U1887 ( .A(n6519), .B(\Variables[0][2][1]_wire ), .C(n6678), 
        .D(\Variables[1][2][1]_wire ), .Z(n6893) );
    GTECH_AOI222 U1888 ( .A(\Variables[2][2][0]_wire ), .B(n6677), .C(
        \Variables[4][2][0]_wire ), .D(n6673), .E(\Variables[3][2][0]_wire ), 
        .F(n6676), .Z(n6894) );
    GTECH_AOI22 U1889 ( .A(n6519), .B(\Variables[0][2][0]_wire ), .C(n6678), 
        .D(\Variables[1][2][0]_wire ), .Z(n6895) );
    GTECH_AOI222 U1890 ( .A(\Variables[2][1][3]_wire ), .B(n6677), .C(
        \Variables[4][1][3]_wire ), .D(n6673), .E(\Variables[3][1][3]_wire ), 
        .F(n6676), .Z(n6896) );
    GTECH_AOI22 U1891 ( .A(n6519), .B(\Variables[0][1][3]_wire ), .C(n6678), 
        .D(\Variables[1][1][3]_wire ), .Z(n6897) );
    GTECH_AOI222 U1892 ( .A(\Variables[2][1][2]_wire ), .B(n6677), .C(
        \Variables[4][1][2]_wire ), .D(n6673), .E(\Variables[3][1][2]_wire ), 
        .F(n6676), .Z(n6898) );
    GTECH_AOI22 U1893 ( .A(n6519), .B(\Variables[0][1][2]_wire ), .C(n6678), 
        .D(\Variables[1][1][2]_wire ), .Z(n6899) );
    GTECH_AOI222 U1894 ( .A(\Variables[2][1][1]_wire ), .B(n6677), .C(
        \Variables[4][1][1]_wire ), .D(n6673), .E(\Variables[3][1][1]_wire ), 
        .F(n6676), .Z(n6900) );
    GTECH_AOI22 U1895 ( .A(n6519), .B(\Variables[0][1][1]_wire ), .C(n6678), 
        .D(\Variables[1][1][1]_wire ), .Z(n6901) );
    GTECH_AOI222 U1896 ( .A(\Variables[2][1][0]_wire ), .B(n6677), .C(
        \Variables[4][1][0]_wire ), .D(n6673), .E(\Variables[3][1][0]_wire ), 
        .F(n6676), .Z(n6902) );
    GTECH_AOI22 U1897 ( .A(n6519), .B(\Variables[0][1][0]_wire ), .C(n6678), 
        .D(\Variables[1][1][0]_wire ), .Z(n6903) );
    GTECH_AOI222 U1898 ( .A(\Variables[2][0][3]_wire ), .B(n6677), .C(
        \Variables[4][0][3]_wire ), .D(n6673), .E(\Variables[3][0][3]_wire ), 
        .F(n6676), .Z(n6904) );
    GTECH_AOI22 U1899 ( .A(n6519), .B(\Variables[0][0][3]_wire ), .C(n6678), 
        .D(\Variables[1][0][3]_wire ), .Z(n6905) );
    GTECH_AOI222 U1900 ( .A(\Variables[2][0][2]_wire ), .B(n6677), .C(
        \Variables[4][0][2]_wire ), .D(n6673), .E(\Variables[3][0][2]_wire ), 
        .F(n6676), .Z(n6906) );
    GTECH_AOI22 U1901 ( .A(n6519), .B(\Variables[0][0][2]_wire ), .C(n6678), 
        .D(\Variables[1][0][2]_wire ), .Z(n6907) );
    GTECH_AOI222 U1902 ( .A(\Variables[2][0][1]_wire ), .B(n6677), .C(
        \Variables[4][0][1]_wire ), .D(n6673), .E(\Variables[3][0][1]_wire ), 
        .F(n6676), .Z(n6908) );
    GTECH_AOI22 U1903 ( .A(n6519), .B(\Variables[0][0][1]_wire ), .C(n6678), 
        .D(\Variables[1][0][1]_wire ), .Z(n6909) );
    GTECH_AOI222 U1904 ( .A(\Variables[2][0][0]_wire ), .B(n6677), .C(
        \Variables[4][0][0]_wire ), .D(n6673), .E(\Variables[3][0][0]_wire ), 
        .F(n6676), .Z(n6910) );
    GTECH_AOI22 U1905 ( .A(n6519), .B(\Variables[0][0][0]_wire ), .C(n6678), 
        .D(\Variables[1][0][0]_wire ), .Z(n6911) );
    GTECH_AOI22 U1906 ( .A(n6673), .B(\Variables[4][-8][3]_wire ), .C(n6676), 
        .D(\Variables[3][-8][3]_wire ), .Z(n6792) );
    GTECH_AOI22 U1907 ( .A(n6677), .B(\Variables[2][-8][3]_wire ), .C(n6678), 
        .D(\Variables[1][-8][3]_wire ), .Z(n6791) );
    GTECH_AOI22 U1908 ( .A(n6673), .B(\Variables[4][-8][2]_wire ), .C(n6676), 
        .D(\Variables[3][-8][2]_wire ), .Z(n6831) );
    GTECH_AOI22 U1909 ( .A(n6677), .B(\Variables[2][-8][2]_wire ), .C(n6678), 
        .D(\Variables[1][-8][2]_wire ), .Z(n6830) );
    GTECH_AOI22 U1910 ( .A(n6673), .B(\Variables[4][-8][1]_wire ), .C(n6676), 
        .D(\Variables[3][-8][1]_wire ), .Z(n6837) );
    GTECH_AOI22 U1911 ( .A(n6677), .B(\Variables[2][-8][1]_wire ), .C(n6678), 
        .D(\Variables[1][-8][1]_wire ), .Z(n6836) );
    GTECH_AOI22 U1912 ( .A(n6673), .B(\Variables[4][-8][0]_wire ), .C(n6676), 
        .D(\Variables[3][-8][0]_wire ), .Z(n6843) );
    GTECH_AOI22 U1913 ( .A(n6677), .B(\Variables[2][-8][0]_wire ), .C(n6678), 
        .D(\Variables[1][-8][0]_wire ), .Z(n6842) );
    GTECH_AOI22 U1914 ( .A(n6673), .B(\Variables[4][-7][3]_wire ), .C(n6676), 
        .D(\Variables[3][-7][3]_wire ), .Z(n6787) );
    GTECH_AOI22 U1915 ( .A(n6677), .B(\Variables[2][-7][3]_wire ), .C(n6678), 
        .D(\Variables[1][-7][3]_wire ), .Z(n6786) );
    GTECH_AOI22 U1916 ( .A(n6673), .B(\Variables[4][-7][2]_wire ), .C(n6676), 
        .D(\Variables[3][-7][2]_wire ), .Z(n6829) );
    GTECH_AOI22 U1917 ( .A(n6677), .B(\Variables[2][-7][2]_wire ), .C(n6678), 
        .D(\Variables[1][-7][2]_wire ), .Z(n6828) );
    GTECH_AOI22 U1918 ( .A(n6673), .B(\Variables[4][-7][1]_wire ), .C(n6676), 
        .D(\Variables[3][-7][1]_wire ), .Z(n6835) );
    GTECH_AOI22 U1919 ( .A(n6677), .B(\Variables[2][-7][1]_wire ), .C(n6678), 
        .D(\Variables[1][-7][1]_wire ), .Z(n6834) );
    GTECH_AOI22 U1920 ( .A(n6673), .B(\Variables[4][-7][0]_wire ), .C(n6676), 
        .D(\Variables[3][-7][0]_wire ), .Z(n6841) );
    GTECH_AOI22 U1921 ( .A(n6677), .B(\Variables[2][-7][0]_wire ), .C(n6678), 
        .D(\Variables[1][-7][0]_wire ), .Z(n6840) );
    GTECH_AOI222 U1922 ( .A(\Variables[2][-6][3]_wire ), .B(n6677), .C(
        \Variables[4][-6][3]_wire ), .D(n6673), .E(\Variables[3][-6][3]_wire ), 
        .F(n6676), .Z(n6912) );
    GTECH_AOI22 U1923 ( .A(n6519), .B(\Variables[0][-6][3]_wire ), .C(n6678), 
        .D(\Variables[1][-6][3]_wire ), .Z(n6913) );
    GTECH_AOI222 U1924 ( .A(\Variables[2][-6][2]_wire ), .B(n6677), .C(
        \Variables[4][-6][2]_wire ), .D(n6673), .E(\Variables[3][-6][2]_wire ), 
        .F(n6676), .Z(n6914) );
    GTECH_AOI22 U1925 ( .A(n6519), .B(\Variables[0][-6][2]_wire ), .C(n6678), 
        .D(\Variables[1][-6][2]_wire ), .Z(n6915) );
    GTECH_AOI222 U1926 ( .A(\Variables[2][-6][1]_wire ), .B(n6677), .C(
        \Variables[4][-6][1]_wire ), .D(n6673), .E(\Variables[3][-6][1]_wire ), 
        .F(n6676), .Z(n6916) );
    GTECH_AOI22 U1927 ( .A(n6519), .B(\Variables[0][-6][1]_wire ), .C(n6678), 
        .D(\Variables[1][-6][1]_wire ), .Z(n6917) );
    GTECH_AOI222 U1928 ( .A(\Variables[2][-6][0]_wire ), .B(n6677), .C(
        \Variables[4][-6][0]_wire ), .D(n6673), .E(\Variables[3][-6][0]_wire ), 
        .F(n6676), .Z(n6918) );
    GTECH_AOI22 U1929 ( .A(n6519), .B(\Variables[0][-6][0]_wire ), .C(n6678), 
        .D(\Variables[1][-6][0]_wire ), .Z(n6919) );
    GTECH_AOI222 U1930 ( .A(\Variables[2][-5][3]_wire ), .B(n6677), .C(
        \Variables[4][-5][3]_wire ), .D(n6673), .E(\Variables[3][-5][3]_wire ), 
        .F(n6676), .Z(n6920) );
    GTECH_AOI22 U1931 ( .A(n6519), .B(\Variables[0][-5][3]_wire ), .C(n6678), 
        .D(\Variables[1][-5][3]_wire ), .Z(n6921) );
    GTECH_AOI222 U1932 ( .A(\Variables[2][-5][2]_wire ), .B(n6677), .C(
        \Variables[4][-5][2]_wire ), .D(n6673), .E(\Variables[3][-5][2]_wire ), 
        .F(n6676), .Z(n6922) );
    GTECH_AOI22 U1933 ( .A(n6519), .B(\Variables[0][-5][2]_wire ), .C(n6678), 
        .D(\Variables[1][-5][2]_wire ), .Z(n6923) );
    GTECH_AOI222 U1934 ( .A(\Variables[2][-5][1]_wire ), .B(n6677), .C(
        \Variables[4][-5][1]_wire ), .D(n6673), .E(\Variables[3][-5][1]_wire ), 
        .F(n6676), .Z(n6924) );
    GTECH_AOI22 U1935 ( .A(n6519), .B(\Variables[0][-5][1]_wire ), .C(n6678), 
        .D(\Variables[1][-5][1]_wire ), .Z(n6925) );
    GTECH_AOI222 U1936 ( .A(\Variables[2][-5][0]_wire ), .B(n6677), .C(
        \Variables[4][-5][0]_wire ), .D(n6673), .E(\Variables[3][-5][0]_wire ), 
        .F(n6676), .Z(n6926) );
    GTECH_AOI22 U1937 ( .A(n6519), .B(\Variables[0][-5][0]_wire ), .C(n6678), 
        .D(\Variables[1][-5][0]_wire ), .Z(n6927) );
    GTECH_AOI222 U1938 ( .A(\Variables[2][-4][3]_wire ), .B(n6677), .C(
        \Variables[4][-4][3]_wire ), .D(n6673), .E(\Variables[3][-4][3]_wire ), 
        .F(n6676), .Z(n6928) );
    GTECH_AOI22 U1939 ( .A(n6519), .B(\Variables[0][-4][3]_wire ), .C(n6678), 
        .D(\Variables[1][-4][3]_wire ), .Z(n6929) );
    GTECH_AOI222 U1940 ( .A(\Variables[2][-4][2]_wire ), .B(n6677), .C(
        \Variables[4][-4][2]_wire ), .D(n6673), .E(\Variables[3][-4][2]_wire ), 
        .F(n6676), .Z(n6930) );
    GTECH_AOI22 U1941 ( .A(n6519), .B(\Variables[0][-4][2]_wire ), .C(n6678), 
        .D(\Variables[1][-4][2]_wire ), .Z(n6931) );
    GTECH_AOI222 U1942 ( .A(\Variables[2][-4][1]_wire ), .B(n6677), .C(
        \Variables[4][-4][1]_wire ), .D(n6673), .E(\Variables[3][-4][1]_wire ), 
        .F(n6676), .Z(n6932) );
    GTECH_AOI22 U1943 ( .A(n6519), .B(\Variables[0][-4][1]_wire ), .C(n6678), 
        .D(\Variables[1][-4][1]_wire ), .Z(n6933) );
    GTECH_AOI222 U1944 ( .A(\Variables[2][-4][0]_wire ), .B(n6677), .C(
        \Variables[4][-4][0]_wire ), .D(n6673), .E(\Variables[3][-4][0]_wire ), 
        .F(n6676), .Z(n6934) );
    GTECH_AOI22 U1945 ( .A(n6519), .B(\Variables[0][-4][0]_wire ), .C(n6678), 
        .D(\Variables[1][-4][0]_wire ), .Z(n6935) );
    GTECH_AOI22 U1946 ( .A(n6673), .B(\Variables[4][-3][3]_wire ), .C(n6676), 
        .D(\Variables[3][-3][3]_wire ), .Z(n6782) );
    GTECH_AOI22 U1947 ( .A(n6677), .B(\Variables[2][-3][3]_wire ), .C(n6678), 
        .D(\Variables[1][-3][3]_wire ), .Z(n6781) );
    GTECH_AOI22 U1948 ( .A(n6673), .B(\Variables[4][-3][2]_wire ), .C(n6676), 
        .D(\Variables[3][-3][2]_wire ), .Z(n6827) );
    GTECH_AOI22 U1949 ( .A(n6677), .B(\Variables[2][-3][2]_wire ), .C(n6678), 
        .D(\Variables[1][-3][2]_wire ), .Z(n6826) );
    GTECH_AOI22 U1950 ( .A(n6673), .B(\Variables[4][-3][1]_wire ), .C(n6676), 
        .D(\Variables[3][-3][1]_wire ), .Z(n6833) );
    GTECH_AOI22 U1951 ( .A(n6677), .B(\Variables[2][-3][1]_wire ), .C(n6678), 
        .D(\Variables[1][-3][1]_wire ), .Z(n6832) );
    GTECH_AOI22 U1952 ( .A(n6673), .B(\Variables[4][-3][0]_wire ), .C(n6676), 
        .D(\Variables[3][-3][0]_wire ), .Z(n6839) );
    GTECH_AOI22 U1953 ( .A(n6677), .B(\Variables[2][-3][0]_wire ), .C(n6678), 
        .D(\Variables[1][-3][0]_wire ), .Z(n6838) );
    GTECH_AOI222 U1954 ( .A(\Variables[2][-2][3]_wire ), .B(n6677), .C(
        \Variables[4][-2][3]_wire ), .D(n6673), .E(\Variables[3][-2][3]_wire ), 
        .F(n6676), .Z(n6936) );
    GTECH_AOI22 U1955 ( .A(n6519), .B(\Variables[0][-2][3]_wire ), .C(n6678), 
        .D(\Variables[1][-2][3]_wire ), .Z(n6937) );
    GTECH_AOI222 U1956 ( .A(\Variables[2][-2][2]_wire ), .B(n6677), .C(
        \Variables[4][-2][2]_wire ), .D(n6673), .E(\Variables[3][-2][2]_wire ), 
        .F(n6676), .Z(n6938) );
    GTECH_AOI22 U1957 ( .A(n6519), .B(\Variables[0][-2][2]_wire ), .C(n6678), 
        .D(\Variables[1][-2][2]_wire ), .Z(n6939) );
    GTECH_AOI222 U1958 ( .A(\Variables[2][-2][1]_wire ), .B(n6677), .C(
        \Variables[4][-2][1]_wire ), .D(n6673), .E(\Variables[3][-2][1]_wire ), 
        .F(n6676), .Z(n6940) );
    GTECH_AOI22 U1959 ( .A(n6519), .B(\Variables[0][-2][1]_wire ), .C(n6678), 
        .D(\Variables[1][-2][1]_wire ), .Z(n6941) );
    GTECH_AOI222 U1960 ( .A(\Variables[2][-2][0]_wire ), .B(n6677), .C(
        \Variables[4][-2][0]_wire ), .D(n6673), .E(\Variables[3][-2][0]_wire ), 
        .F(n6676), .Z(n6942) );
    GTECH_AOI22 U1961 ( .A(n6519), .B(\Variables[0][-2][0]_wire ), .C(n6678), 
        .D(\Variables[1][-2][0]_wire ), .Z(n6943) );
    GTECH_AOI222 U1962 ( .A(\Variables[2][-1][3]_wire ), .B(n6677), .C(
        \Variables[4][-1][3]_wire ), .D(n6673), .E(\Variables[3][-1][3]_wire ), 
        .F(n6676), .Z(n6944) );
    GTECH_AOI22 U1963 ( .A(n6519), .B(\Variables[0][-1][3]_wire ), .C(n6678), 
        .D(\Variables[1][-1][3]_wire ), .Z(n6945) );
    GTECH_AOI222 U1964 ( .A(\Variables[2][-1][2]_wire ), .B(n6677), .C(
        \Variables[4][-1][2]_wire ), .D(n6673), .E(\Variables[3][-1][2]_wire ), 
        .F(n6676), .Z(n6946) );
    GTECH_AOI22 U1965 ( .A(n6519), .B(\Variables[0][-1][2]_wire ), .C(n6678), 
        .D(\Variables[1][-1][2]_wire ), .Z(n6947) );
    GTECH_AOI222 U1966 ( .A(\Variables[2][-1][1]_wire ), .B(n6677), .C(
        \Variables[4][-1][1]_wire ), .D(n6673), .E(\Variables[3][-1][1]_wire ), 
        .F(n6676), .Z(n6948) );
    GTECH_AOI22 U1967 ( .A(n6678), .B(\Variables[1][-1][1]_wire ), .C(n6519), 
        .D(\Variables[0][-1][1]_wire ), .Z(n6949) );
    GTECH_AOI222 U1968 ( .A(\Variables[2][-1][0]_wire ), .B(n6677), .C(
        \Variables[4][-1][0]_wire ), .D(n6673), .E(\Variables[3][-1][0]_wire ), 
        .F(n6676), .Z(n6950) );
    GTECH_AOI22 U1969 ( .A(n6519), .B(\Variables[0][-1][0]_wire ), .C(n6678), 
        .D(\Variables[1][-1][0]_wire ), .Z(n6951) );
    GTECH_AOI222 U1970 ( .A(n6725), .B(\Variables[2][7][3]_wire ), .C(n6721), 
        .D(\Variables[4][7][3]_wire ), .E(n6724), .F(\Variables[3][7][3]_wire 
        ), .Z(n6952) );
    GTECH_AOI22 U1971 ( .A(\Variables[0][7][3]_wire ), .B(n6727), .C(
        \Variables[1][7][3]_wire ), .D(n6726), .Z(n6953) );
    GTECH_AOI222 U1972 ( .A(n6725), .B(\Variables[2][6][3]_wire ), .C(n6721), 
        .D(\Variables[4][6][3]_wire ), .E(n6724), .F(\Variables[3][6][3]_wire 
        ), .Z(n6954) );
    GTECH_AOI22 U1973 ( .A(\Variables[0][6][3]_wire ), .B(n6727), .C(
        \Variables[1][6][3]_wire ), .D(n6726), .Z(n6955) );
    GTECH_AOI222 U1974 ( .A(n6725), .B(\Variables[2][5][3]_wire ), .C(n6721), 
        .D(\Variables[4][5][3]_wire ), .E(n6724), .F(\Variables[3][5][3]_wire 
        ), .Z(n6956) );
    GTECH_AOI22 U1975 ( .A(\Variables[0][5][3]_wire ), .B(n6727), .C(
        \Variables[1][5][3]_wire ), .D(n6726), .Z(n6957) );
    GTECH_AOI222 U1976 ( .A(n6725), .B(\Variables[2][4][3]_wire ), .C(n6721), 
        .D(\Variables[4][4][3]_wire ), .E(n6724), .F(\Variables[3][4][3]_wire 
        ), .Z(n6958) );
    GTECH_AOI22 U1977 ( .A(\Variables[0][4][3]_wire ), .B(n6727), .C(
        \Variables[1][4][3]_wire ), .D(n6726), .Z(n6959) );
    GTECH_AOI222 U1978 ( .A(n6725), .B(\Variables[2][3][3]_wire ), .C(n6721), 
        .D(\Variables[4][3][3]_wire ), .E(n6724), .F(\Variables[3][3][3]_wire 
        ), .Z(n6960) );
    GTECH_AOI22 U1979 ( .A(\Variables[0][3][3]_wire ), .B(n6727), .C(
        \Variables[1][3][3]_wire ), .D(n6726), .Z(n6961) );
    GTECH_AOI222 U1980 ( .A(n6725), .B(\Variables[2][2][3]_wire ), .C(n6721), 
        .D(\Variables[4][2][3]_wire ), .E(n6724), .F(\Variables[3][2][3]_wire 
        ), .Z(n6962) );
    GTECH_AOI22 U1981 ( .A(\Variables[0][2][3]_wire ), .B(n6727), .C(
        \Variables[1][2][3]_wire ), .D(n6726), .Z(n6963) );
    GTECH_AOI222 U1982 ( .A(n6725), .B(\Variables[2][1][3]_wire ), .C(n6721), 
        .D(\Variables[4][1][3]_wire ), .E(n6724), .F(\Variables[3][1][3]_wire 
        ), .Z(n6964) );
    GTECH_AOI22 U1983 ( .A(\Variables[0][1][3]_wire ), .B(n6727), .C(
        \Variables[1][1][3]_wire ), .D(n6726), .Z(n6965) );
    GTECH_AOI222 U1984 ( .A(n6725), .B(\Variables[2][0][3]_wire ), .C(n6721), 
        .D(\Variables[4][0][3]_wire ), .E(n6724), .F(\Variables[3][0][3]_wire 
        ), .Z(n6966) );
    GTECH_AOI22 U1985 ( .A(\Variables[0][0][3]_wire ), .B(n6727), .C(
        \Variables[1][0][3]_wire ), .D(n6726), .Z(n6967) );
    GTECH_AOI222 U1986 ( .A(n6725), .B(\Variables[2][-1][3]_wire ), .C(n6721), 
        .D(\Variables[4][-1][3]_wire ), .E(n6724), .F(
        \Variables[3][-1][3]_wire ), .Z(n6968) );
    GTECH_AOI22 U1987 ( .A(\Variables[0][-1][3]_wire ), .B(n6727), .C(
        \Variables[1][-1][3]_wire ), .D(n6726), .Z(n6969) );
    GTECH_AOI222 U1988 ( .A(n6725), .B(\Variables[2][-2][3]_wire ), .C(n6721), 
        .D(\Variables[4][-2][3]_wire ), .E(n6724), .F(
        \Variables[3][-2][3]_wire ), .Z(n6970) );
    GTECH_AOI22 U1989 ( .A(\Variables[0][-2][3]_wire ), .B(n6727), .C(
        \Variables[1][-2][3]_wire ), .D(n6726), .Z(n6971) );
    GTECH_AOI222 U1990 ( .A(n6725), .B(\Variables[2][-3][3]_wire ), .C(n6721), 
        .D(\Variables[4][-3][3]_wire ), .E(n6724), .F(
        \Variables[3][-3][3]_wire ), .Z(n6972) );
    GTECH_AOI22 U1991 ( .A(\Variables[1][-3][3]_wire ), .B(n6726), .C(
        \Variables[0][-3][3]_wire ), .D(n6727), .Z(n6973) );
    GTECH_AOI222 U1992 ( .A(n6725), .B(\Variables[2][-4][3]_wire ), .C(n6721), 
        .D(\Variables[4][-4][3]_wire ), .E(n6724), .F(
        \Variables[3][-4][3]_wire ), .Z(n6974) );
    GTECH_AOI22 U1993 ( .A(\Variables[0][-4][3]_wire ), .B(n6727), .C(
        \Variables[1][-4][3]_wire ), .D(n6726), .Z(n6975) );
    GTECH_AOI222 U1994 ( .A(n6725), .B(\Variables[2][-5][3]_wire ), .C(n6721), 
        .D(\Variables[4][-5][3]_wire ), .E(n6724), .F(
        \Variables[3][-5][3]_wire ), .Z(n6976) );
    GTECH_AOI22 U1995 ( .A(\Variables[0][-5][3]_wire ), .B(n6727), .C(
        \Variables[1][-5][3]_wire ), .D(n6726), .Z(n6977) );
    GTECH_AOI222 U1996 ( .A(n6725), .B(\Variables[2][-6][3]_wire ), .C(n6721), 
        .D(\Variables[4][-6][3]_wire ), .E(n6724), .F(
        \Variables[3][-6][3]_wire ), .Z(n6978) );
    GTECH_AOI22 U1997 ( .A(\Variables[0][-6][3]_wire ), .B(n6727), .C(
        \Variables[1][-6][3]_wire ), .D(n6726), .Z(n6979) );
    GTECH_AOI222 U1998 ( .A(n6725), .B(\Variables[2][-7][3]_wire ), .C(n6721), 
        .D(\Variables[4][-7][3]_wire ), .E(n6724), .F(
        \Variables[3][-7][3]_wire ), .Z(n6980) );
    GTECH_AOI22 U1999 ( .A(\Variables[1][-7][3]_wire ), .B(n6726), .C(
        \Variables[0][-7][3]_wire ), .D(n6727), .Z(n6981) );
    GTECH_AOI222 U2000 ( .A(n6725), .B(\Variables[2][-8][3]_wire ), .C(n6721), 
        .D(\Variables[4][-8][3]_wire ), .E(n6724), .F(
        \Variables[3][-8][3]_wire ), .Z(n6982) );
    GTECH_AOI22 U2001 ( .A(\Variables[1][-8][3]_wire ), .B(n6726), .C(
        \Variables[0][-8][3]_wire ), .D(n6727), .Z(n6983) );
    GTECH_OA22 U2002 ( .A(n6984), .B(n6730), .C(n6985), .D(n6728), .Z(n6547)
         );
    GTECH_AOI2N2 U2003 ( .A(n6986), .B(n6734), .C(n6987), .D(n6732), .Z(n6546)
         );
    GTECH_AOI2N2 U2004 ( .A(n6988), .B(n6737), .C(n6989), .D(n6736), .Z(n6545)
         );
    GTECH_AOI2N2 U2005 ( .A(n6990), .B(n6739), .C(n6991), .D(n6738), .Z(n6544)
         );
    GTECH_AOI2N2 U2006 ( .A(n6992), .B(n6742), .C(n6993), .D(n6741), .Z(n6543)
         );
    GTECH_AOI2N2 U2007 ( .A(n6994), .B(n6744), .C(n6995), .D(n6743), .Z(n6542)
         );
    GTECH_AOI2N2 U2008 ( .A(n6996), .B(n6997), .C(n6998), .D(n6746), .Z(n6541)
         );
    GTECH_OA22 U2009 ( .A(n6999), .B(n6749), .C(n7000), .D(n6748), .Z(n6540)
         );
    GTECH_AOI222 U2010 ( .A(n6725), .B(\Variables[2][7][2]_wire ), .C(n6721), 
        .D(\Variables[4][7][2]_wire ), .E(n6724), .F(\Variables[3][7][2]_wire 
        ), .Z(n7001) );
    GTECH_AOI22 U2011 ( .A(\Variables[0][7][2]_wire ), .B(n6727), .C(
        \Variables[1][7][2]_wire ), .D(n6726), .Z(n7002) );
    GTECH_AOI222 U2012 ( .A(n6725), .B(\Variables[2][6][2]_wire ), .C(n6721), 
        .D(\Variables[4][6][2]_wire ), .E(n6724), .F(\Variables[3][6][2]_wire 
        ), .Z(n7003) );
    GTECH_AOI22 U2013 ( .A(\Variables[0][6][2]_wire ), .B(n6727), .C(
        \Variables[1][6][2]_wire ), .D(n6726), .Z(n7004) );
    GTECH_AOI222 U2014 ( .A(n6725), .B(\Variables[2][5][2]_wire ), .C(n6721), 
        .D(\Variables[4][5][2]_wire ), .E(n6724), .F(\Variables[3][5][2]_wire 
        ), .Z(n7005) );
    GTECH_AOI22 U2015 ( .A(\Variables[0][5][2]_wire ), .B(n6727), .C(
        \Variables[1][5][2]_wire ), .D(n6726), .Z(n7006) );
    GTECH_AOI222 U2016 ( .A(n6725), .B(\Variables[2][4][2]_wire ), .C(n6721), 
        .D(\Variables[4][4][2]_wire ), .E(n6724), .F(\Variables[3][4][2]_wire 
        ), .Z(n7007) );
    GTECH_AOI22 U2017 ( .A(\Variables[0][4][2]_wire ), .B(n6727), .C(
        \Variables[1][4][2]_wire ), .D(n6726), .Z(n7008) );
    GTECH_AOI222 U2018 ( .A(n6725), .B(\Variables[2][3][2]_wire ), .C(n6721), 
        .D(\Variables[4][3][2]_wire ), .E(n6724), .F(\Variables[3][3][2]_wire 
        ), .Z(n7009) );
    GTECH_AOI22 U2019 ( .A(\Variables[0][3][2]_wire ), .B(n6727), .C(
        \Variables[1][3][2]_wire ), .D(n6726), .Z(n7010) );
    GTECH_AOI222 U2020 ( .A(n6725), .B(\Variables[2][2][2]_wire ), .C(n6721), 
        .D(\Variables[4][2][2]_wire ), .E(n6724), .F(\Variables[3][2][2]_wire 
        ), .Z(n7011) );
    GTECH_AOI22 U2021 ( .A(\Variables[0][2][2]_wire ), .B(n6727), .C(
        \Variables[1][2][2]_wire ), .D(n6726), .Z(n7012) );
    GTECH_AOI222 U2022 ( .A(n6725), .B(\Variables[2][1][2]_wire ), .C(n6721), 
        .D(\Variables[4][1][2]_wire ), .E(n6724), .F(\Variables[3][1][2]_wire 
        ), .Z(n7013) );
    GTECH_AOI22 U2023 ( .A(\Variables[0][1][2]_wire ), .B(n6727), .C(
        \Variables[1][1][2]_wire ), .D(n6726), .Z(n7014) );
    GTECH_AOI222 U2024 ( .A(n6725), .B(\Variables[2][0][2]_wire ), .C(n6721), 
        .D(\Variables[4][0][2]_wire ), .E(n6724), .F(\Variables[3][0][2]_wire 
        ), .Z(n7015) );
    GTECH_AOI22 U2025 ( .A(\Variables[0][0][2]_wire ), .B(n6727), .C(
        \Variables[1][0][2]_wire ), .D(n6726), .Z(n7016) );
    GTECH_AOI222 U2026 ( .A(n6725), .B(\Variables[2][-1][2]_wire ), .C(n6721), 
        .D(\Variables[4][-1][2]_wire ), .E(n6724), .F(
        \Variables[3][-1][2]_wire ), .Z(n7017) );
    GTECH_AOI22 U2027 ( .A(\Variables[0][-1][2]_wire ), .B(n6727), .C(
        \Variables[1][-1][2]_wire ), .D(n6726), .Z(n7018) );
    GTECH_AOI222 U2028 ( .A(n6725), .B(\Variables[2][-2][2]_wire ), .C(n6721), 
        .D(\Variables[4][-2][2]_wire ), .E(n6724), .F(
        \Variables[3][-2][2]_wire ), .Z(n7019) );
    GTECH_AOI22 U2029 ( .A(\Variables[0][-2][2]_wire ), .B(n6727), .C(
        \Variables[1][-2][2]_wire ), .D(n6726), .Z(n7020) );
    GTECH_AOI222 U2030 ( .A(n6725), .B(\Variables[2][-3][2]_wire ), .C(n6721), 
        .D(\Variables[4][-3][2]_wire ), .E(n6724), .F(
        \Variables[3][-3][2]_wire ), .Z(n7021) );
    GTECH_AOI22 U2031 ( .A(\Variables[1][-3][2]_wire ), .B(n6726), .C(
        \Variables[0][-3][2]_wire ), .D(n6727), .Z(n7022) );
    GTECH_AOI222 U2032 ( .A(n6725), .B(\Variables[2][-4][2]_wire ), .C(n6721), 
        .D(\Variables[4][-4][2]_wire ), .E(n6724), .F(
        \Variables[3][-4][2]_wire ), .Z(n7023) );
    GTECH_AOI22 U2033 ( .A(\Variables[0][-4][2]_wire ), .B(n6727), .C(
        \Variables[1][-4][2]_wire ), .D(n6726), .Z(n7024) );
    GTECH_AOI222 U2034 ( .A(n6725), .B(\Variables[2][-5][2]_wire ), .C(n6721), 
        .D(\Variables[4][-5][2]_wire ), .E(n6724), .F(
        \Variables[3][-5][2]_wire ), .Z(n7025) );
    GTECH_AOI22 U2035 ( .A(\Variables[0][-5][2]_wire ), .B(n6727), .C(
        \Variables[1][-5][2]_wire ), .D(n6726), .Z(n7026) );
    GTECH_AOI222 U2036 ( .A(n6725), .B(\Variables[2][-6][2]_wire ), .C(n6721), 
        .D(\Variables[4][-6][2]_wire ), .E(n6724), .F(
        \Variables[3][-6][2]_wire ), .Z(n7027) );
    GTECH_AOI22 U2037 ( .A(\Variables[0][-6][2]_wire ), .B(n6727), .C(
        \Variables[1][-6][2]_wire ), .D(n6726), .Z(n7028) );
    GTECH_AOI222 U2038 ( .A(n6725), .B(\Variables[2][-7][2]_wire ), .C(n6721), 
        .D(\Variables[4][-7][2]_wire ), .E(n6724), .F(
        \Variables[3][-7][2]_wire ), .Z(n7029) );
    GTECH_AOI22 U2039 ( .A(\Variables[1][-7][2]_wire ), .B(n6726), .C(
        \Variables[0][-7][2]_wire ), .D(n6727), .Z(n7030) );
    GTECH_AOI222 U2040 ( .A(n6725), .B(\Variables[2][-8][2]_wire ), .C(n6721), 
        .D(\Variables[4][-8][2]_wire ), .E(n6724), .F(
        \Variables[3][-8][2]_wire ), .Z(n7031) );
    GTECH_AOI22 U2041 ( .A(\Variables[1][-8][2]_wire ), .B(n6726), .C(
        \Variables[0][-8][2]_wire ), .D(n6727), .Z(n7032) );
    GTECH_OA22 U2042 ( .A(n7033), .B(n6730), .C(n7034), .D(n6728), .Z(n6555)
         );
    GTECH_AOI2N2 U2043 ( .A(n7035), .B(n6734), .C(n7036), .D(n6732), .Z(n6554)
         );
    GTECH_AOI2N2 U2044 ( .A(n7037), .B(n6737), .C(n7038), .D(n6736), .Z(n6553)
         );
    GTECH_AOI2N2 U2045 ( .A(n7039), .B(n6739), .C(n7040), .D(n6738), .Z(n6552)
         );
    GTECH_AOI2N2 U2046 ( .A(n7041), .B(n6742), .C(n7042), .D(n6741), .Z(n6551)
         );
    GTECH_AOI2N2 U2047 ( .A(n7043), .B(n6744), .C(n7044), .D(n6743), .Z(n6550)
         );
    GTECH_AOI2N2 U2048 ( .A(n7045), .B(n6997), .C(n7046), .D(n6746), .Z(n6549)
         );
    GTECH_OA22 U2049 ( .A(n7047), .B(n6749), .C(n7048), .D(n6748), .Z(n6548)
         );
    GTECH_AOI222 U2050 ( .A(n6725), .B(\Variables[2][7][1]_wire ), .C(n6721), 
        .D(\Variables[4][7][1]_wire ), .E(n6724), .F(\Variables[3][7][1]_wire 
        ), .Z(n7049) );
    GTECH_AOI22 U2051 ( .A(\Variables[0][7][1]_wire ), .B(n6727), .C(
        \Variables[1][7][1]_wire ), .D(n6726), .Z(n7050) );
    GTECH_AOI222 U2052 ( .A(n6725), .B(\Variables[2][6][1]_wire ), .C(n6721), 
        .D(\Variables[4][6][1]_wire ), .E(n6724), .F(\Variables[3][6][1]_wire 
        ), .Z(n7051) );
    GTECH_AOI22 U2053 ( .A(\Variables[0][6][1]_wire ), .B(n6727), .C(
        \Variables[1][6][1]_wire ), .D(n6726), .Z(n7052) );
    GTECH_AOI222 U2054 ( .A(n6725), .B(\Variables[2][5][1]_wire ), .C(n6721), 
        .D(\Variables[4][5][1]_wire ), .E(n6724), .F(\Variables[3][5][1]_wire 
        ), .Z(n7053) );
    GTECH_AOI22 U2055 ( .A(\Variables[0][5][1]_wire ), .B(n6727), .C(
        \Variables[1][5][1]_wire ), .D(n6726), .Z(n7054) );
    GTECH_AOI222 U2056 ( .A(n6725), .B(\Variables[2][4][1]_wire ), .C(n6721), 
        .D(\Variables[4][4][1]_wire ), .E(n6724), .F(\Variables[3][4][1]_wire 
        ), .Z(n7055) );
    GTECH_AOI22 U2057 ( .A(\Variables[0][4][1]_wire ), .B(n6727), .C(
        \Variables[1][4][1]_wire ), .D(n6726), .Z(n7056) );
    GTECH_AOI222 U2058 ( .A(n6725), .B(\Variables[2][3][1]_wire ), .C(n6721), 
        .D(\Variables[4][3][1]_wire ), .E(n6724), .F(\Variables[3][3][1]_wire 
        ), .Z(n7057) );
    GTECH_AOI22 U2059 ( .A(\Variables[0][3][1]_wire ), .B(n6727), .C(
        \Variables[1][3][1]_wire ), .D(n6726), .Z(n7058) );
    GTECH_AOI222 U2060 ( .A(n6725), .B(\Variables[2][2][1]_wire ), .C(n6721), 
        .D(\Variables[4][2][1]_wire ), .E(n6724), .F(\Variables[3][2][1]_wire 
        ), .Z(n7059) );
    GTECH_AOI22 U2061 ( .A(\Variables[0][2][1]_wire ), .B(n6727), .C(
        \Variables[1][2][1]_wire ), .D(n6726), .Z(n7060) );
    GTECH_AOI222 U2062 ( .A(n6725), .B(\Variables[2][1][1]_wire ), .C(n6721), 
        .D(\Variables[4][1][1]_wire ), .E(n6724), .F(\Variables[3][1][1]_wire 
        ), .Z(n7061) );
    GTECH_AOI22 U2063 ( .A(\Variables[0][1][1]_wire ), .B(n6727), .C(
        \Variables[1][1][1]_wire ), .D(n6726), .Z(n7062) );
    GTECH_AOI222 U2064 ( .A(n6725), .B(\Variables[2][0][1]_wire ), .C(n6721), 
        .D(\Variables[4][0][1]_wire ), .E(n6724), .F(\Variables[3][0][1]_wire 
        ), .Z(n7063) );
    GTECH_AOI22 U2065 ( .A(\Variables[0][0][1]_wire ), .B(n6727), .C(
        \Variables[1][0][1]_wire ), .D(n6726), .Z(n7064) );
    GTECH_AOI222 U2066 ( .A(n6725), .B(\Variables[2][-1][1]_wire ), .C(n6721), 
        .D(\Variables[4][-1][1]_wire ), .E(n6724), .F(
        \Variables[3][-1][1]_wire ), .Z(n7065) );
    GTECH_AOI22 U2067 ( .A(\Variables[1][-1][1]_wire ), .B(n6726), .C(
        \Variables[0][-1][1]_wire ), .D(n6727), .Z(n7066) );
    GTECH_AOI222 U2068 ( .A(n6725), .B(\Variables[2][-2][1]_wire ), .C(n6721), 
        .D(\Variables[4][-2][1]_wire ), .E(n6724), .F(
        \Variables[3][-2][1]_wire ), .Z(n7067) );
    GTECH_AOI22 U2069 ( .A(\Variables[0][-2][1]_wire ), .B(n6727), .C(
        \Variables[1][-2][1]_wire ), .D(n6726), .Z(n7068) );
    GTECH_AOI222 U2070 ( .A(n6725), .B(\Variables[2][-3][1]_wire ), .C(n6721), 
        .D(\Variables[4][-3][1]_wire ), .E(n6724), .F(
        \Variables[3][-3][1]_wire ), .Z(n7069) );
    GTECH_AOI22 U2071 ( .A(\Variables[1][-3][1]_wire ), .B(n6726), .C(
        \Variables[0][-3][1]_wire ), .D(n6727), .Z(n7070) );
    GTECH_AOI222 U2072 ( .A(n6725), .B(\Variables[2][-4][1]_wire ), .C(n6721), 
        .D(\Variables[4][-4][1]_wire ), .E(n6724), .F(
        \Variables[3][-4][1]_wire ), .Z(n7071) );
    GTECH_AOI22 U2073 ( .A(\Variables[0][-4][1]_wire ), .B(n6727), .C(
        \Variables[1][-4][1]_wire ), .D(n6726), .Z(n7072) );
    GTECH_AOI222 U2074 ( .A(n6725), .B(\Variables[2][-5][1]_wire ), .C(n6721), 
        .D(\Variables[4][-5][1]_wire ), .E(n6724), .F(
        \Variables[3][-5][1]_wire ), .Z(n7073) );
    GTECH_AOI22 U2075 ( .A(\Variables[0][-5][1]_wire ), .B(n6727), .C(
        \Variables[1][-5][1]_wire ), .D(n6726), .Z(n7074) );
    GTECH_AOI222 U2076 ( .A(n6725), .B(\Variables[2][-6][1]_wire ), .C(n6721), 
        .D(\Variables[4][-6][1]_wire ), .E(n6724), .F(
        \Variables[3][-6][1]_wire ), .Z(n7075) );
    GTECH_AOI22 U2077 ( .A(\Variables[0][-6][1]_wire ), .B(n6727), .C(
        \Variables[1][-6][1]_wire ), .D(n6726), .Z(n7076) );
    GTECH_AOI222 U2078 ( .A(n6725), .B(\Variables[2][-7][1]_wire ), .C(n6721), 
        .D(\Variables[4][-7][1]_wire ), .E(n6724), .F(
        \Variables[3][-7][1]_wire ), .Z(n7077) );
    GTECH_AOI22 U2079 ( .A(\Variables[1][-7][1]_wire ), .B(n6726), .C(
        \Variables[0][-7][1]_wire ), .D(n6727), .Z(n7078) );
    GTECH_AOI222 U2080 ( .A(n6725), .B(\Variables[2][-8][1]_wire ), .C(n6721), 
        .D(\Variables[4][-8][1]_wire ), .E(n6724), .F(
        \Variables[3][-8][1]_wire ), .Z(n7079) );
    GTECH_AOI22 U2081 ( .A(\Variables[1][-8][1]_wire ), .B(n6726), .C(
        \Variables[0][-8][1]_wire ), .D(n6727), .Z(n7080) );
    GTECH_OA22 U2082 ( .A(n7081), .B(n6730), .C(n7082), .D(n6728), .Z(n6563)
         );
    GTECH_AOI2N2 U2083 ( .A(n7083), .B(n6734), .C(n7084), .D(n6732), .Z(n6562)
         );
    GTECH_AOI2N2 U2084 ( .A(n7085), .B(n6737), .C(n7086), .D(n6736), .Z(n6561)
         );
    GTECH_AOI2N2 U2085 ( .A(n7087), .B(n6739), .C(n7088), .D(n6738), .Z(n6560)
         );
    GTECH_AOI2N2 U2086 ( .A(n7089), .B(n6742), .C(n7090), .D(n6741), .Z(n6559)
         );
    GTECH_AOI2N2 U2087 ( .A(n7091), .B(n6744), .C(n7092), .D(n6743), .Z(n6558)
         );
    GTECH_AOI2N2 U2088 ( .A(n7093), .B(n6997), .C(n7094), .D(n6746), .Z(n6557)
         );
    GTECH_OA22 U2089 ( .A(n7095), .B(n6749), .C(n7096), .D(n6748), .Z(n6556)
         );
    GTECH_AOI222 U2090 ( .A(n6725), .B(\Variables[2][7][0]_wire ), .C(n6721), 
        .D(\Variables[4][7][0]_wire ), .E(n6724), .F(\Variables[3][7][0]_wire 
        ), .Z(n7097) );
    GTECH_AOI22 U2091 ( .A(\Variables[0][7][0]_wire ), .B(n6727), .C(
        \Variables[1][7][0]_wire ), .D(n6726), .Z(n7098) );
    GTECH_AOI222 U2092 ( .A(n6725), .B(\Variables[2][6][0]_wire ), .C(n6721), 
        .D(\Variables[4][6][0]_wire ), .E(n6724), .F(\Variables[3][6][0]_wire 
        ), .Z(n7099) );
    GTECH_AOI22 U2093 ( .A(\Variables[1][6][0]_wire ), .B(n6726), .C(
        \Variables[0][6][0]_wire ), .D(n6727), .Z(n7100) );
    GTECH_AOI222 U2094 ( .A(n6725), .B(\Variables[2][5][0]_wire ), .C(n6721), 
        .D(\Variables[4][5][0]_wire ), .E(n6724), .F(\Variables[3][5][0]_wire 
        ), .Z(n7101) );
    GTECH_AOI22 U2095 ( .A(\Variables[0][5][0]_wire ), .B(n6727), .C(
        \Variables[1][5][0]_wire ), .D(n6726), .Z(n7102) );
    GTECH_AOI222 U2096 ( .A(n6725), .B(\Variables[2][4][0]_wire ), .C(n6721), 
        .D(\Variables[4][4][0]_wire ), .E(n6724), .F(\Variables[3][4][0]_wire 
        ), .Z(n7103) );
    GTECH_AOI22 U2097 ( .A(\Variables[0][4][0]_wire ), .B(n6727), .C(
        \Variables[1][4][0]_wire ), .D(n6726), .Z(n7104) );
    GTECH_AOI222 U2098 ( .A(n6725), .B(\Variables[2][3][0]_wire ), .C(n6721), 
        .D(\Variables[4][3][0]_wire ), .E(n6724), .F(\Variables[3][3][0]_wire 
        ), .Z(n7105) );
    GTECH_AOI22 U2099 ( .A(\Variables[0][3][0]_wire ), .B(n6727), .C(
        \Variables[1][3][0]_wire ), .D(n6726), .Z(n7106) );
    GTECH_AOI222 U2100 ( .A(n6725), .B(\Variables[2][2][0]_wire ), .C(n6721), 
        .D(\Variables[4][2][0]_wire ), .E(n6724), .F(\Variables[3][2][0]_wire 
        ), .Z(n7107) );
    GTECH_AOI22 U2101 ( .A(\Variables[0][2][0]_wire ), .B(n6727), .C(
        \Variables[1][2][0]_wire ), .D(n6726), .Z(n7108) );
    GTECH_AOI222 U2102 ( .A(n6725), .B(\Variables[2][1][0]_wire ), .C(n6721), 
        .D(\Variables[4][1][0]_wire ), .E(n6724), .F(\Variables[3][1][0]_wire 
        ), .Z(n7109) );
    GTECH_AOI22 U2103 ( .A(\Variables[0][1][0]_wire ), .B(n6727), .C(
        \Variables[1][1][0]_wire ), .D(n6726), .Z(n7110) );
    GTECH_AOI222 U2104 ( .A(n6725), .B(\Variables[2][0][0]_wire ), .C(n6721), 
        .D(\Variables[4][0][0]_wire ), .E(n6724), .F(\Variables[3][0][0]_wire 
        ), .Z(n7111) );
    GTECH_AOI22 U2105 ( .A(\Variables[0][0][0]_wire ), .B(n6727), .C(
        \Variables[1][0][0]_wire ), .D(n6726), .Z(n7112) );
    GTECH_AOI222 U2106 ( .A(n6725), .B(\Variables[2][-1][0]_wire ), .C(n6721), 
        .D(\Variables[4][-1][0]_wire ), .E(n6724), .F(
        \Variables[3][-1][0]_wire ), .Z(n7113) );
    GTECH_AOI22 U2107 ( .A(\Variables[0][-1][0]_wire ), .B(n6727), .C(
        \Variables[1][-1][0]_wire ), .D(n6726), .Z(n7114) );
    GTECH_AOI222 U2108 ( .A(n6725), .B(\Variables[2][-2][0]_wire ), .C(n6721), 
        .D(\Variables[4][-2][0]_wire ), .E(n6724), .F(
        \Variables[3][-2][0]_wire ), .Z(n7115) );
    GTECH_AOI22 U2109 ( .A(\Variables[0][-2][0]_wire ), .B(n6727), .C(
        \Variables[1][-2][0]_wire ), .D(n6726), .Z(n7116) );
    GTECH_AOI222 U2110 ( .A(n6725), .B(\Variables[2][-3][0]_wire ), .C(n6721), 
        .D(\Variables[4][-3][0]_wire ), .E(n6724), .F(
        \Variables[3][-3][0]_wire ), .Z(n7117) );
    GTECH_AOI22 U2111 ( .A(\Variables[1][-3][0]_wire ), .B(n6726), .C(
        \Variables[0][-3][0]_wire ), .D(n6727), .Z(n7118) );
    GTECH_AOI222 U2112 ( .A(n6725), .B(\Variables[2][-4][0]_wire ), .C(n6721), 
        .D(\Variables[4][-4][0]_wire ), .E(n6724), .F(
        \Variables[3][-4][0]_wire ), .Z(n7119) );
    GTECH_AOI22 U2113 ( .A(\Variables[0][-4][0]_wire ), .B(n6727), .C(
        \Variables[1][-4][0]_wire ), .D(n6726), .Z(n7120) );
    GTECH_AOI222 U2114 ( .A(n6725), .B(\Variables[2][-5][0]_wire ), .C(n6721), 
        .D(\Variables[4][-5][0]_wire ), .E(n6724), .F(
        \Variables[3][-5][0]_wire ), .Z(n7121) );
    GTECH_AOI22 U2115 ( .A(\Variables[0][-5][0]_wire ), .B(n6727), .C(
        \Variables[1][-5][0]_wire ), .D(n6726), .Z(n7122) );
    GTECH_AOI222 U2116 ( .A(n6725), .B(\Variables[2][-6][0]_wire ), .C(n6721), 
        .D(\Variables[4][-6][0]_wire ), .E(n6724), .F(
        \Variables[3][-6][0]_wire ), .Z(n7123) );
    GTECH_AOI22 U2117 ( .A(\Variables[0][-6][0]_wire ), .B(n6727), .C(
        \Variables[1][-6][0]_wire ), .D(n6726), .Z(n7124) );
    GTECH_AOI222 U2118 ( .A(n6725), .B(\Variables[2][-7][0]_wire ), .C(n6721), 
        .D(\Variables[4][-7][0]_wire ), .E(n6724), .F(
        \Variables[3][-7][0]_wire ), .Z(n7125) );
    GTECH_AOI22 U2119 ( .A(\Variables[1][-7][0]_wire ), .B(n6726), .C(
        \Variables[0][-7][0]_wire ), .D(n6727), .Z(n7126) );
    GTECH_AOI222 U2120 ( .A(n6725), .B(\Variables[2][-8][0]_wire ), .C(n6721), 
        .D(\Variables[4][-8][0]_wire ), .E(n6724), .F(
        \Variables[3][-8][0]_wire ), .Z(n7127) );
    GTECH_AOI22 U2121 ( .A(\Variables[1][-8][0]_wire ), .B(n6726), .C(
        \Variables[0][-8][0]_wire ), .D(n6727), .Z(n7128) );
    GTECH_OA22 U2122 ( .A(n7129), .B(n6730), .C(n7130), .D(n6728), .Z(n6571)
         );
    GTECH_AOI2N2 U2123 ( .A(n7131), .B(n6734), .C(n7132), .D(n6732), .Z(n6570)
         );
    GTECH_AOI2N2 U2124 ( .A(n7133), .B(n6737), .C(n7134), .D(n6736), .Z(n6569)
         );
    GTECH_AOI2N2 U2125 ( .A(n7135), .B(n6739), .C(n7136), .D(n6738), .Z(n6568)
         );
    GTECH_AOI2N2 U2126 ( .A(n7137), .B(n6742), .C(n7138), .D(n6741), .Z(n6567)
         );
    GTECH_AOI2N2 U2127 ( .A(n7139), .B(n6744), .C(n7140), .D(n6743), .Z(n6566)
         );
    GTECH_OA22 U2128 ( .A(n7141), .B(n6747), .C(n7142), .D(n6746), .Z(n6565)
         );
    GTECH_OA22 U2129 ( .A(n7143), .B(n6749), .C(n7144), .D(n6748), .Z(n6564)
         );
    GTECH_AND2 U2130 ( .A(n6728), .B(n6745), .Z(n6751) );
    GTECH_OA22 U2131 ( .A(n6984), .B(n6757), .C(n6985), .D(n6755), .Z(n6579)
         );
    GTECH_AOI2N2 U2132 ( .A(n6986), .B(n6761), .C(n6987), .D(n6760), .Z(n6578)
         );
    GTECH_AOI2N2 U2133 ( .A(n6988), .B(n6765), .C(n6989), .D(n6763), .Z(n6577)
         );
    GTECH_AOI2N2 U2134 ( .A(n6990), .B(n6767), .C(n6991), .D(n6766), .Z(n6576)
         );
    GTECH_AOI2N2 U2135 ( .A(n6992), .B(n6770), .C(n6993), .D(n6769), .Z(n6575)
         );
    GTECH_AOI2N2 U2136 ( .A(n6994), .B(n6773), .C(n6995), .D(n6772), .Z(n6574)
         );
    GTECH_OA22 U2137 ( .A(n7145), .B(n7146), .C(n6998), .D(n6774), .Z(n6573)
         );
    GTECH_OA22 U2138 ( .A(n6999), .B(n6777), .C(n7000), .D(n6776), .Z(n6572)
         );
    GTECH_OA22 U2139 ( .A(n7033), .B(n6757), .C(n7034), .D(n6755), .Z(n6587)
         );
    GTECH_AOI2N2 U2140 ( .A(n7035), .B(n6761), .C(n7036), .D(n6760), .Z(n6586)
         );
    GTECH_AOI2N2 U2141 ( .A(n7037), .B(n6765), .C(n7038), .D(n6763), .Z(n6585)
         );
    GTECH_AOI2N2 U2142 ( .A(n7039), .B(n6767), .C(n7040), .D(n6766), .Z(n6584)
         );
    GTECH_AOI2N2 U2143 ( .A(n7041), .B(n6770), .C(n7042), .D(n6769), .Z(n6583)
         );
    GTECH_AOI2N2 U2144 ( .A(n7043), .B(n6773), .C(n7044), .D(n6772), .Z(n6582)
         );
    GTECH_OA22 U2145 ( .A(n7147), .B(n7146), .C(n7046), .D(n6774), .Z(n6581)
         );
    GTECH_OA22 U2146 ( .A(n7047), .B(n6777), .C(n7048), .D(n6776), .Z(n6580)
         );
    GTECH_OA22 U2147 ( .A(n7081), .B(n6757), .C(n7082), .D(n6755), .Z(n6595)
         );
    GTECH_AOI2N2 U2148 ( .A(n7083), .B(n6761), .C(n7084), .D(n6760), .Z(n6594)
         );
    GTECH_AOI2N2 U2149 ( .A(n7085), .B(n6765), .C(n7086), .D(n6763), .Z(n6593)
         );
    GTECH_AOI2N2 U2150 ( .A(n7087), .B(n6767), .C(n7088), .D(n6766), .Z(n6592)
         );
    GTECH_AOI2N2 U2151 ( .A(n7089), .B(n6770), .C(n7090), .D(n6769), .Z(n6591)
         );
    GTECH_AOI2N2 U2152 ( .A(n7091), .B(n6773), .C(n7092), .D(n6772), .Z(n6590)
         );
    GTECH_AOI2N2 U2153 ( .A(n7093), .B(n6775), .C(n7094), .D(n6774), .Z(n6589)
         );
    GTECH_OA22 U2154 ( .A(n7095), .B(n6777), .C(n7096), .D(n6776), .Z(n6588)
         );
    GTECH_OA22 U2155 ( .A(n7130), .B(n6755), .C(n7129), .D(n6757), .Z(n6603)
         );
    GTECH_AOI2N2 U2156 ( .A(n7131), .B(n6761), .C(n7132), .D(n6760), .Z(n6602)
         );
    GTECH_AOI2N2 U2157 ( .A(n7133), .B(n6765), .C(n7134), .D(n6763), .Z(n6601)
         );
    GTECH_AOI2N2 U2158 ( .A(n7135), .B(n6767), .C(n7136), .D(n6766), .Z(n6600)
         );
    GTECH_AOI2N2 U2159 ( .A(n7137), .B(n6770), .C(n7138), .D(n6769), .Z(n6599)
         );
    GTECH_AOI2N2 U2160 ( .A(n7139), .B(n6773), .C(n7140), .D(n6772), .Z(n6598)
         );
    GTECH_OA22 U2161 ( .A(n7142), .B(n6774), .C(n7141), .D(n7146), .Z(n6597)
         );
    GTECH_OA22 U2162 ( .A(n7144), .B(n6776), .C(n7143), .D(n6777), .Z(n6596)
         );
    GTECH_OA22 U2163 ( .A(n7340), .B(n7148), .C(n7337), .D(n7149), .Z(n6483)
         );
    GTECH_OA22 U2164 ( .A(n7148), .B(n7339), .C(n6318), .D(n7338), .Z(n6478)
         );
    GTECH_OA22 U2165 ( .A(ReturnJump), .B(n6480), .C(n7149), .D(n7336), .Z(
        n6477) );
    GTECH_OA22 U2166 ( .A(n7151), .B(n7152), .C(n7153), .D(n6783), .Z(n7150)
         );
    GTECH_AOI2N2 U2167 ( .A(n7155), .B(n6795), .C(n7156), .D(n6793), .Z(n7154)
         );
    GTECH_AOI22 U2168 ( .A(n7158), .B(n6797), .C(n7159), .D(n6799), .Z(n7157)
         );
    GTECH_AOI22 U2169 ( .A(n7161), .B(n6800), .C(n7162), .D(n6801), .Z(n7160)
         );
    GTECH_AOI22 U2170 ( .A(n7164), .B(n6802), .C(n7165), .D(n6803), .Z(n7163)
         );
    GTECH_AOI2N2 U2171 ( .A(n7167), .B(n6804), .C(n7168), .D(n6806), .Z(n7166)
         );
    GTECH_AOI22 U2172 ( .A(n7170), .B(n6807), .C(n7171), .D(n6808), .Z(n7169)
         );
    GTECH_AOI22 U2173 ( .A(n7173), .B(n6809), .C(n7174), .D(n6810), .Z(n7172)
         );
    GTECH_AOI222 U2174 ( .A(n6449), .B(n6619), .C(\product1846[5] ), .D(n6448), 
        .E(n6812), .F(n6617), .Z(n7175) );
    GTECH_AOI222 U2175 ( .A(\Lower[3] ), .B(n6845), .C(n6818), .D(\Upper[3] ), 
        .E(n6332), .F(\Lower[2] ), .Z(n7176) );
    GTECH_OA21 U2176 ( .A(n6663), .B(n7178), .C(n6651), .Z(n7177) );
    GTECH_OA21 U2177 ( .A(n6667), .B(n6844), .C(n7180), .Z(n7179) );
    GTECH_AOI2N2 U2178 ( .A(n7182), .B(n6820), .C(n7153), .D(n6819), .Z(n7181)
         );
    GTECH_AOI2N2 U2179 ( .A(n7155), .B(n6330), .C(n7156), .D(n6821), .Z(n7183)
         );
    GTECH_AOI22 U2180 ( .A(n7158), .B(n6822), .C(n7159), .D(n6812), .Z(n7184)
         );
    GTECH_AOI22 U2181 ( .A(n7161), .B(n6332), .C(n6845), .D(n7162), .Z(n7185)
         );
    GTECH_AOI22 U2182 ( .A(n7164), .B(n6449), .C(n7165), .D(n6448), .Z(n7186)
         );
    GTECH_AOI2N2 U2183 ( .A(n7167), .B(n6635), .C(n7168), .D(n6823), .Z(n7187)
         );
    GTECH_AOI22 U2184 ( .A(n7170), .B(n6824), .C(n7171), .D(n6618), .Z(n7188)
         );
    GTECH_AOI22 U2185 ( .A(n7173), .B(n6818), .C(n7174), .D(n6431), .Z(n7189)
         );
    GTECH_AOI222 U2186 ( .A(n6669), .B(n7191), .C(\TableSelect[3] ), .D(n6778), 
        .E(n6811), .F(n7192), .Z(n7190) );
    GTECH_AOI222 U2187 ( .A(n6487), .B(n7194), .C(MemoryReadValue[3]), .D(
        n7195), .E(n6486), .F(\NextInstruction[PARAMETER][3] ), .Z(n7193) );
    GTECH_OA22 U2188 ( .A(n7197), .B(n7152), .C(n7198), .D(n6783), .Z(n7196)
         );
    GTECH_OA22 U2189 ( .A(n7200), .B(n7201), .C(n7202), .D(n6793), .Z(n7199)
         );
    GTECH_AOI22 U2190 ( .A(n7204), .B(n6797), .C(n7205), .D(n6799), .Z(n7203)
         );
    GTECH_AOI22 U2191 ( .A(n7207), .B(n6800), .C(n7208), .D(n6801), .Z(n7206)
         );
    GTECH_AOI22 U2192 ( .A(n7210), .B(n6802), .C(n7211), .D(n6803), .Z(n7209)
         );
    GTECH_AOI2N2 U2193 ( .A(n7213), .B(n6804), .C(n7214), .D(n6806), .Z(n7212)
         );
    GTECH_AOI22 U2194 ( .A(n7216), .B(n6807), .C(n7217), .D(n6808), .Z(n7215)
         );
    GTECH_AOI22 U2195 ( .A(n7219), .B(n6809), .C(n7220), .D(n6810), .Z(n7218)
         );
    GTECH_AOI222 U2196 ( .A(n6449), .B(n6621), .C(\product1846[4] ), .D(n6448), 
        .E(n6812), .F(n6620), .Z(n7221) );
    GTECH_AOI222 U2197 ( .A(\Lower[3] ), .B(n6845), .C(n6818), .D(\Upper[2] ), 
        .E(n6332), .F(\Lower[1] ), .Z(n7222) );
    GTECH_OA22 U2198 ( .A(n7198), .B(n6819), .C(n7197), .D(n7224), .Z(n7223)
         );
    GTECH_OA22 U2199 ( .A(n7200), .B(n7226), .C(n7202), .D(n6821), .Z(n7225)
         );
    GTECH_AOI22 U2200 ( .A(n7204), .B(n6822), .C(n7205), .D(n6812), .Z(n7227)
         );
    GTECH_AOI22 U2201 ( .A(n7207), .B(n6332), .C(n6845), .D(n7208), .Z(n7228)
         );
    GTECH_AOI22 U2202 ( .A(n7210), .B(n6449), .C(n7211), .D(n6448), .Z(n7229)
         );
    GTECH_AOI2N2 U2203 ( .A(n7213), .B(n6635), .C(n7214), .D(n6823), .Z(n7230)
         );
    GTECH_AOI22 U2204 ( .A(n7216), .B(n6824), .C(n7217), .D(n6618), .Z(n7231)
         );
    GTECH_AOI22 U2205 ( .A(n7219), .B(n6818), .C(n7220), .D(n6431), .Z(n7232)
         );
    GTECH_AOI222 U2206 ( .A(n6669), .B(n7234), .C(n6778), .D(\gt_236/AEQB[2] ), 
        .E(n6811), .F(n7235), .Z(n7233) );
    GTECH_AOI222 U2207 ( .A(n6487), .B(n7237), .C(MemoryReadValue[2]), .D(
        n7195), .E(n6486), .F(\NextInstruction[PARAMETER][2] ), .Z(n7236) );
    GTECH_AOI2N2 U2208 ( .A(n7239), .B(n6788), .C(n7240), .D(n6783), .Z(n7238)
         );
    GTECH_OA22 U2209 ( .A(n7242), .B(n6793), .C(n7243), .D(n7201), .Z(n7241)
         );
    GTECH_AOI22 U2210 ( .A(n7245), .B(n6797), .C(n7246), .D(n6799), .Z(n7244)
         );
    GTECH_AOI22 U2211 ( .A(n7248), .B(n6801), .C(n7249), .D(n6800), .Z(n7247)
         );
    GTECH_AOI22 U2212 ( .A(n7251), .B(n6802), .C(n7252), .D(n6803), .Z(n7250)
         );
    GTECH_AOI2N2 U2213 ( .A(n7254), .B(n6804), .C(n7255), .D(n6806), .Z(n7253)
         );
    GTECH_AOI22 U2214 ( .A(n7257), .B(n6808), .C(n7258), .D(n6807), .Z(n7256)
         );
    GTECH_AOI22 U2215 ( .A(n7260), .B(n6809), .C(n7261), .D(n6810), .Z(n7259)
         );
    GTECH_AOI222 U2216 ( .A(n6623), .B(n6449), .C(\product1846[3] ), .D(n6448), 
        .E(n6812), .F(n6622), .Z(n7262) );
    GTECH_AOI222 U2217 ( .A(\Lower[2] ), .B(n6845), .C(n6818), .D(\Upper[1] ), 
        .E(n6332), .F(\Lower[0] ), .Z(n7263) );
    GTECH_AOI2N2 U2218 ( .A(n7239), .B(n6820), .C(n7240), .D(n6819), .Z(n7264)
         );
    GTECH_OA22 U2219 ( .A(n7243), .B(n7226), .C(n7242), .D(n6821), .Z(n7265)
         );
    GTECH_AOI22 U2220 ( .A(n7245), .B(n6822), .C(n7246), .D(n6812), .Z(n7266)
         );
    GTECH_AOI22 U2221 ( .A(n7249), .B(n6332), .C(n6845), .D(n7248), .Z(n7267)
         );
    GTECH_AOI22 U2222 ( .A(n7251), .B(n6449), .C(n7252), .D(n6448), .Z(n7268)
         );
    GTECH_AOI2N2 U2223 ( .A(n7254), .B(n6635), .C(n7255), .D(n6823), .Z(n7269)
         );
    GTECH_AOI22 U2224 ( .A(n7258), .B(n6824), .C(n7257), .D(n6618), .Z(n7270)
         );
    GTECH_AOI22 U2225 ( .A(n7260), .B(n6818), .C(n7261), .D(n6431), .Z(n7271)
         );
    GTECH_AOI222 U2226 ( .A(n6669), .B(n7273), .C(n6778), .D(\TableSelect[1] ), 
        .E(n6811), .F(n7274), .Z(n7272) );
    GTECH_AOI222 U2227 ( .A(n6487), .B(n7276), .C(MemoryReadValue[1]), .D(
        n7195), .E(n6486), .F(\NextInstruction[PARAMETER][1] ), .Z(n7275) );
    GTECH_OA22 U2228 ( .A(n7278), .B(n6783), .C(n7279), .D(n7152), .Z(n7277)
         );
    GTECH_AOI2N2 U2229 ( .A(n7281), .B(n6795), .C(n7282), .D(n6793), .Z(n7280)
         );
    GTECH_AOI22 U2230 ( .A(n7284), .B(n6797), .C(n7285), .D(n6799), .Z(n7283)
         );
    GTECH_AOI22 U2231 ( .A(n7287), .B(n6800), .C(n7288), .D(n6801), .Z(n7286)
         );
    GTECH_AOI22 U2232 ( .A(n7290), .B(n6802), .C(n7291), .D(n6803), .Z(n7289)
         );
    GTECH_AOI2N2 U2233 ( .A(n7293), .B(n6804), .C(n7294), .D(n6806), .Z(n7292)
         );
    GTECH_AOI22 U2234 ( .A(n7296), .B(n6807), .C(n7297), .D(n6808), .Z(n7295)
         );
    GTECH_AOI22 U2235 ( .A(n7299), .B(n6809), .C(n7300), .D(n6810), .Z(n7298)
         );
    GTECH_AOI222 U2236 ( .A(n6449), .B(n6625), .C(\product1846[2] ), .D(n6448), 
        .E(n6812), .F(n6624), .Z(n7301) );
    GTECH_AOI22 U2237 ( .A(\Upper[0] ), .B(n6818), .C(n6845), .D(\Lower[1] ), 
        .Z(n7302) );
    GTECH_OA22 U2238 ( .A(n7278), .B(n6819), .C(n7279), .D(n7224), .Z(n7303)
         );
    GTECH_AOI2N2 U2239 ( .A(n7281), .B(n6330), .C(n7282), .D(n6821), .Z(n7304)
         );
    GTECH_AOI22 U2240 ( .A(n7284), .B(n6822), .C(n7285), .D(n6812), .Z(n7305)
         );
    GTECH_AOI22 U2241 ( .A(n7287), .B(n6332), .C(n6845), .D(n7288), .Z(n7306)
         );
    GTECH_AOI22 U2242 ( .A(n7290), .B(n6449), .C(n7291), .D(n6448), .Z(n7307)
         );
    GTECH_AOI2N2 U2243 ( .A(n7293), .B(n6635), .C(n7294), .D(n6823), .Z(n7308)
         );
    GTECH_AOI22 U2244 ( .A(n7296), .B(n6824), .C(n7297), .D(n6618), .Z(n7309)
         );
    GTECH_AOI22 U2245 ( .A(n7299), .B(n6818), .C(n7300), .D(n6431), .Z(n7310)
         );
    GTECH_AOI222 U2246 ( .A(n6669), .B(n7312), .C(n6778), .D(\TableSelect[0] ), 
        .E(n6811), .F(n7313), .Z(n7311) );
    GTECH_AOI222 U2247 ( .A(n6487), .B(n7315), .C(MemoryReadValue[0]), .D(
        n7195), .E(n6486), .F(\NextInstruction[PARAMETER][0] ), .Z(n7314) );
    GTECH_AND2 U2248 ( .A(n7316), .B(n6652), .Z(n6629) );
    GTECH_OAI21 U2249 ( .A(n6626), .B(n6651), .C(n7317), .Z(n6327) );
    GTECH_OAI21 U2250 ( .A(\NextInstruction[PARAMETER][2] ), .B(n6630), .C(
        n6427), .Z(n7318) );
    GTECH_OA21 U2251 ( .A(n6633), .B(n7318), .C(n6627), .Z(n6334) );
    GTECH_OR_NOT U2252 ( .A(n6701), .B(n6696), .Z(n6637) );
    GTECH_NAND2 U2253 ( .A(n6702), .B(n6696), .Z(n6638) );
    GTECH_OR_NOT U2254 ( .A(n6685), .B(n6702), .Z(n6639) );
    GTECH_NOT U2255 ( .A(IRQInProcess), .Z(n6473) );
    GTECH_NOT U2256 ( .A(n6519), .Z(n6713) );
    GTECH_NOT U2257 ( .A(n6328), .Z(n6471) );
    GTECH_NOT U2258 ( .A(ResetStarted), .Z(n6322) );
    GTECH_NOT U2259 ( .A(ReturnJump), .Z(n6481) );
    GTECH_NOT U2260 ( .A(n6669), .Z(n6844) );
    GTECH_NOT U2261 ( .A(n6819), .Z(n6616) );
    GTECH_NOT U2262 ( .A(n6427), .Z(n6845) );
    GTECH_NOT U2263 ( .A(n_660), .Z(n6320) );
    GTECH_AND_NOT U2264 ( .A(\Upper[3] ), .B(n6336), .Z(n7319) );
    GTECH_AND2 U2265 ( .A(\NextInstruction[PARAMETER][3] ), .B(\Upper[2] ), 
        .Z(n6817) );
    GTECH_AND2 U2266 ( .A(\Upper[1] ), .B(\NextInstruction[PARAMETER][3] ), 
        .Z(n6814) );
    GTECH_NOT U2267 ( .A(n6659), .Z(n6665) );
    GTECH_AND2 U2268 ( .A(\Upper[0] ), .B(\NextInstruction[PARAMETER][3] ), 
        .Z(n6614) );
    GTECH_NOT U2269 ( .A(n6475), .Z(n6649) );
    GTECH_OR3 U2270 ( .A(\IRQ[3] ), .B(\IRQ[4] ), .C(n6649), .Z(n6647) );
    GTECH_OR3 U2271 ( .A(n6649), .B(\IRQ[3] ), .C(n6320), .Z(n6648) );
    GTECH_NAND5 U2272 ( .A(IRQCLKEnable), .B(n_399), .C(n_398), .D(n_397), .E(
        n6847), .Z(n6319) );
    GTECH_NAND3 U2273 ( .A(n_660), .B(n6325), .C(\IRQ[1] ), .Z(n6324) );
    GTECH_OAI21 U2274 ( .A(n6812), .B(n6822), .C(n6329), .Z(n6459) );
    GTECH_NAND3 U2275 ( .A(\NextInstruction[INSTRUCTION][2] ), .B(n6650), .C(
        n6660), .Z(n6457) );
    GTECH_NAND3 U2276 ( .A(n6328), .B(n6845), .C(n6662), .Z(n6458) );
    GTECH_NAND3 U2277 ( .A(n6628), .B(n6655), .C(n6489), .Z(n6666) );
    GTECH_NAND2 U2278 ( .A(n7179), .B(n7177), .Z(n7195) );
    GTECH_OAI21 U2279 ( .A(\NextInstruction[PARAMETER][0] ), .B(n6655), .C(
        n6489), .Z(n7320) );
    GTECH_NAND5 U2280 ( .A(n7320), .B(n6665), .C(n6328), .D(n6669), .E(
        \NextInstruction[PARAMETER][3] ), .Z(n6670) );
    GTECH_NAND2 U2281 ( .A(n6848), .B(n6849), .Z(n7155) );
    GTECH_AOI22 U2282 ( .A(n7155), .B(n6679), .C(\Lower[3] ), .D(n6680), .Z(
        n6399) );
    GTECH_AND2 U2283 ( .A(n6850), .B(n6851), .Z(n7200) );
    GTECH_OA22 U2284 ( .A(n6681), .B(n6453), .C(n7200), .D(n7321), .Z(n6400)
         );
    GTECH_AND2 U2285 ( .A(n6853), .B(n6852), .Z(n7243) );
    GTECH_AOI2N2 U2286 ( .A(n6680), .B(\Lower[1] ), .C(n7243), .D(n7321), .Z(
        n6401) );
    GTECH_NAND2 U2287 ( .A(n6855), .B(n6854), .Z(n7281) );
    GTECH_AOI22 U2288 ( .A(n7281), .B(n6679), .C(n6680), .D(\Lower[0] ), .Z(
        n6402) );
    GTECH_NAND2 U2289 ( .A(n6857), .B(n6856), .Z(n7158) );
    GTECH_AOI22 U2290 ( .A(n7158), .B(n6683), .C(\Lower[3] ), .D(n7322), .Z(
        n6395) );
    GTECH_NAND2 U2291 ( .A(n6859), .B(n6858), .Z(n7204) );
    GTECH_AOI22 U2292 ( .A(n7204), .B(n6683), .C(\Lower[2] ), .D(n7322), .Z(
        n6396) );
    GTECH_NAND2 U2293 ( .A(n6861), .B(n6860), .Z(n7245) );
    GTECH_AOI2N2 U2294 ( .A(n7245), .B(n6683), .C(n6455), .D(n6684), .Z(n6397)
         );
    GTECH_NAND2 U2295 ( .A(n6863), .B(n6862), .Z(n7284) );
    GTECH_AOI22 U2296 ( .A(n7284), .B(n6683), .C(\Lower[0] ), .D(n7322), .Z(
        n6398) );
    GTECH_NAND2 U2297 ( .A(n6864), .B(n6865), .Z(n7159) );
    GTECH_AOI22 U2298 ( .A(\Lower[3] ), .B(n6688), .C(n7159), .D(n6687), .Z(
        n6391) );
    GTECH_NAND2 U2299 ( .A(n6866), .B(n6867), .Z(n7205) );
    GTECH_AOI22 U2300 ( .A(\Lower[2] ), .B(n6688), .C(n7205), .D(n6687), .Z(
        n6392) );
    GTECH_NAND2 U2301 ( .A(n6869), .B(n6868), .Z(n7246) );
    GTECH_AOI22 U2302 ( .A(\Lower[1] ), .B(n6688), .C(n7246), .D(n6687), .Z(
        n6393) );
    GTECH_NAND2 U2303 ( .A(n6871), .B(n6870), .Z(n7285) );
    GTECH_AOI22 U2304 ( .A(\Lower[0] ), .B(n6688), .C(n7285), .D(n6687), .Z(
        n6394) );
    GTECH_NAND2 U2305 ( .A(n6873), .B(n6872), .Z(n7161) );
    GTECH_AOI22 U2306 ( .A(n7161), .B(n6689), .C(\Lower[3] ), .D(n6690), .Z(
        n6387) );
    GTECH_NAND2 U2307 ( .A(n6875), .B(n6874), .Z(n7207) );
    GTECH_AOI22 U2308 ( .A(n7207), .B(n6689), .C(\Lower[2] ), .D(n6690), .Z(
        n6388) );
    GTECH_NAND2 U2309 ( .A(n6877), .B(n6876), .Z(n7249) );
    GTECH_AOI22 U2310 ( .A(n7249), .B(n6689), .C(\Lower[1] ), .D(n6690), .Z(
        n6389) );
    GTECH_NAND2 U2311 ( .A(n6879), .B(n6878), .Z(n7287) );
    GTECH_AOI22 U2312 ( .A(n7287), .B(n6689), .C(\Lower[0] ), .D(n6690), .Z(
        n6390) );
    GTECH_NAND2 U2313 ( .A(n6880), .B(n6881), .Z(n7162) );
    GTECH_AOI2N2 U2314 ( .A(n7162), .B(n6692), .C(n6450), .D(n6693), .Z(n6383)
         );
    GTECH_NAND2 U2315 ( .A(n6882), .B(n6883), .Z(n7208) );
    GTECH_AOI2N2 U2316 ( .A(n7208), .B(n6692), .C(n6453), .D(n6693), .Z(n6384)
         );
    GTECH_NAND2 U2317 ( .A(n6885), .B(n6884), .Z(n7248) );
    GTECH_AOI2N2 U2318 ( .A(n7248), .B(n6692), .C(n6455), .D(n6693), .Z(n6385)
         );
    GTECH_NAND2 U2319 ( .A(n6887), .B(n6886), .Z(n7288) );
    GTECH_AOI2N2 U2320 ( .A(n7288), .B(n6692), .C(n6456), .D(n6693), .Z(n6386)
         );
    GTECH_NAND2 U2321 ( .A(n6889), .B(n6888), .Z(n7164) );
    GTECH_AOI22 U2322 ( .A(n7164), .B(n6694), .C(\Lower[3] ), .D(n7323), .Z(
        n6379) );
    GTECH_NAND2 U2323 ( .A(n6891), .B(n6890), .Z(n7210) );
    GTECH_AOI22 U2324 ( .A(n7210), .B(n6694), .C(\Lower[2] ), .D(n7323), .Z(
        n6380) );
    GTECH_NAND2 U2325 ( .A(n6893), .B(n6892), .Z(n7251) );
    GTECH_AOI2N2 U2326 ( .A(n7251), .B(n6694), .C(n6455), .D(n6695), .Z(n6381)
         );
    GTECH_NAND2 U2327 ( .A(n6895), .B(n6894), .Z(n7290) );
    GTECH_AOI22 U2328 ( .A(n7290), .B(n6694), .C(\Lower[0] ), .D(n7323), .Z(
        n6382) );
    GTECH_NAND2 U2329 ( .A(n6896), .B(n6897), .Z(n7165) );
    GTECH_AOI22 U2330 ( .A(\Lower[3] ), .B(n6698), .C(n7165), .D(n6697), .Z(
        n6375) );
    GTECH_NAND2 U2331 ( .A(n6898), .B(n6899), .Z(n7211) );
    GTECH_AOI22 U2332 ( .A(\Lower[2] ), .B(n6698), .C(n7211), .D(n6697), .Z(
        n6376) );
    GTECH_NAND2 U2333 ( .A(n6901), .B(n6900), .Z(n7252) );
    GTECH_AOI22 U2334 ( .A(\Lower[1] ), .B(n6698), .C(n7252), .D(n6697), .Z(
        n6377) );
    GTECH_NAND2 U2335 ( .A(n6903), .B(n6902), .Z(n7291) );
    GTECH_AOI22 U2336 ( .A(\Lower[0] ), .B(n6698), .C(n7291), .D(n6697), .Z(
        n6378) );
    GTECH_NAND2 U2337 ( .A(n6905), .B(n6904), .Z(n7167) );
    GTECH_AOI22 U2338 ( .A(\Lower[3] ), .B(n6700), .C(n7167), .D(n6699), .Z(
        n6371) );
    GTECH_NAND2 U2339 ( .A(n6907), .B(n6906), .Z(n7213) );
    GTECH_AOI22 U2340 ( .A(\Lower[2] ), .B(n6700), .C(n7213), .D(n6699), .Z(
        n6372) );
    GTECH_NAND2 U2341 ( .A(n6909), .B(n6908), .Z(n7254) );
    GTECH_AOI22 U2342 ( .A(\Lower[1] ), .B(n6700), .C(n7254), .D(n6699), .Z(
        n6373) );
    GTECH_NAND2 U2343 ( .A(n6911), .B(n6910), .Z(n7293) );
    GTECH_AOI22 U2344 ( .A(\Lower[0] ), .B(n6700), .C(n7293), .D(n6699), .Z(
        n6374) );
    GTECH_NAND2 U2345 ( .A(n6912), .B(n6913), .Z(n7174) );
    GTECH_AOI2N2 U2346 ( .A(n7174), .B(n6703), .C(n6450), .D(n6704), .Z(n6345)
         );
    GTECH_NAND2 U2347 ( .A(n6914), .B(n6915), .Z(n7220) );
    GTECH_AOI2N2 U2348 ( .A(n7220), .B(n6703), .C(n6453), .D(n6704), .Z(n6348)
         );
    GTECH_NAND2 U2349 ( .A(n6917), .B(n6916), .Z(n7261) );
    GTECH_AOI2N2 U2350 ( .A(n7261), .B(n6703), .C(n6455), .D(n6704), .Z(n6349)
         );
    GTECH_NAND2 U2351 ( .A(n6918), .B(n6919), .Z(n7300) );
    GTECH_AOI2N2 U2352 ( .A(n7300), .B(n6703), .C(n6456), .D(n6704), .Z(n6350)
         );
    GTECH_NAND2 U2353 ( .A(n6921), .B(n6920), .Z(n7173) );
    GTECH_AOI22 U2354 ( .A(n7173), .B(n6705), .C(\Lower[3] ), .D(n6706), .Z(
        n6351) );
    GTECH_NAND2 U2355 ( .A(n6923), .B(n6922), .Z(n7219) );
    GTECH_AOI22 U2356 ( .A(n7219), .B(n6705), .C(\Lower[2] ), .D(n6706), .Z(
        n6352) );
    GTECH_NAND2 U2357 ( .A(n6925), .B(n6924), .Z(n7260) );
    GTECH_AOI22 U2358 ( .A(n7260), .B(n6705), .C(\Lower[1] ), .D(n6706), .Z(
        n6353) );
    GTECH_NAND2 U2359 ( .A(n6927), .B(n6926), .Z(n7299) );
    GTECH_AOI22 U2360 ( .A(n7299), .B(n6705), .C(\Lower[0] ), .D(n6706), .Z(
        n6354) );
    GTECH_NAND2 U2361 ( .A(n6928), .B(n6929), .Z(n7171) );
    GTECH_AOI2N2 U2362 ( .A(n7171), .B(n6707), .C(n6450), .D(n6708), .Z(n6355)
         );
    GTECH_NAND2 U2363 ( .A(n6930), .B(n6931), .Z(n7217) );
    GTECH_AOI2N2 U2364 ( .A(n7217), .B(n6707), .C(n6453), .D(n6708), .Z(n6356)
         );
    GTECH_NAND2 U2365 ( .A(n6933), .B(n6932), .Z(n7257) );
    GTECH_AOI2N2 U2366 ( .A(n7257), .B(n6707), .C(n6455), .D(n6708), .Z(n6357)
         );
    GTECH_NAND2 U2367 ( .A(n6934), .B(n6935), .Z(n7297) );
    GTECH_AOI2N2 U2368 ( .A(n7297), .B(n6707), .C(n6456), .D(n6708), .Z(n6358)
         );
    GTECH_NAND2 U2369 ( .A(n6937), .B(n6936), .Z(n7170) );
    GTECH_AOI22 U2370 ( .A(n7170), .B(n6709), .C(\Lower[3] ), .D(n6710), .Z(
        n6363) );
    GTECH_NAND2 U2371 ( .A(n6939), .B(n6938), .Z(n7216) );
    GTECH_AOI22 U2372 ( .A(n7216), .B(n6709), .C(\Lower[2] ), .D(n6710), .Z(
        n6364) );
    GTECH_NAND2 U2373 ( .A(n6941), .B(n6940), .Z(n7258) );
    GTECH_AOI22 U2374 ( .A(n7258), .B(n6709), .C(\Lower[1] ), .D(n6710), .Z(
        n6365) );
    GTECH_NAND2 U2375 ( .A(n6943), .B(n6942), .Z(n7296) );
    GTECH_AOI22 U2376 ( .A(n7296), .B(n6709), .C(\Lower[0] ), .D(n6710), .Z(
        n6366) );
    GTECH_AND2 U2377 ( .A(n6945), .B(n6944), .Z(n7168) );
    GTECH_AOI2N2 U2378 ( .A(\Lower[3] ), .B(n6712), .C(n7168), .D(n6711), .Z(
        n6367) );
    GTECH_AND2 U2379 ( .A(n6947), .B(n6946), .Z(n7214) );
    GTECH_AOI2N2 U2380 ( .A(\Lower[2] ), .B(n6712), .C(n7214), .D(n6711), .Z(
        n6368) );
    GTECH_AND2 U2381 ( .A(n6949), .B(n6948), .Z(n7255) );
    GTECH_AOI2N2 U2382 ( .A(\Lower[1] ), .B(n6712), .C(n7255), .D(n6711), .Z(
        n6369) );
    GTECH_AND2 U2383 ( .A(n6951), .B(n6950), .Z(n7294) );
    GTECH_AOI2N2 U2384 ( .A(\Lower[0] ), .B(n6712), .C(n7294), .D(n6711), .Z(
        n6370) );
    GTECH_NAND3 U2385 ( .A(n6652), .B(n6322), .C(
        \NextInstruction[PARAMETER][3] ), .Z(n6452) );
    GTECH_NAND3 U2386 ( .A(n6652), .B(n6322), .C(
        \NextInstruction[PARAMETER][2] ), .Z(n6454) );
    GTECH_OAI21 U2387 ( .A(\TableSelect[0] ), .B(\TableSelect[1] ), .C(
        \gt_236/AEQB[2] ), .Z(n6316) );
    GTECH_AND2 U2388 ( .A(n6982), .B(n6983), .Z(n6999) );
    GTECH_AND2 U2389 ( .A(n6980), .B(n6981), .Z(n7000) );
    GTECH_AND2 U2390 ( .A(n6978), .B(n6979), .Z(n7145) );
    GTECH_AND2 U2391 ( .A(n6976), .B(n6977), .Z(n6998) );
    GTECH_NAND2 U2392 ( .A(n6974), .B(n6975), .Z(n6994) );
    GTECH_AND2 U2393 ( .A(n6972), .B(n6973), .Z(n6995) );
    GTECH_NAND2 U2394 ( .A(n6970), .B(n6971), .Z(n6992) );
    GTECH_AND2 U2395 ( .A(n6968), .B(n6969), .Z(n6993) );
    GTECH_NAND2 U2396 ( .A(n6966), .B(n6967), .Z(n6990) );
    GTECH_AND2 U2397 ( .A(n6964), .B(n6965), .Z(n6991) );
    GTECH_NAND2 U2398 ( .A(n6962), .B(n6963), .Z(n6988) );
    GTECH_AND2 U2399 ( .A(n6960), .B(n6961), .Z(n6989) );
    GTECH_NAND2 U2400 ( .A(n6958), .B(n6959), .Z(n6986) );
    GTECH_AND2 U2401 ( .A(n6956), .B(n6957), .Z(n6987) );
    GTECH_AND2 U2402 ( .A(n6954), .B(n6955), .Z(n6984) );
    GTECH_AND2 U2403 ( .A(n6952), .B(n6953), .Z(n6985) );
    GTECH_AND2 U2404 ( .A(n7031), .B(n7032), .Z(n7047) );
    GTECH_AND2 U2405 ( .A(n7029), .B(n7030), .Z(n7048) );
    GTECH_AND2 U2406 ( .A(n7027), .B(n7028), .Z(n7147) );
    GTECH_AND2 U2407 ( .A(n7025), .B(n7026), .Z(n7046) );
    GTECH_NAND2 U2408 ( .A(n7023), .B(n7024), .Z(n7043) );
    GTECH_AND2 U2409 ( .A(n7021), .B(n7022), .Z(n7044) );
    GTECH_NAND2 U2410 ( .A(n7019), .B(n7020), .Z(n7041) );
    GTECH_AND2 U2411 ( .A(n7017), .B(n7018), .Z(n7042) );
    GTECH_NAND2 U2412 ( .A(n7015), .B(n7016), .Z(n7039) );
    GTECH_AND2 U2413 ( .A(n7013), .B(n7014), .Z(n7040) );
    GTECH_NAND2 U2414 ( .A(n7011), .B(n7012), .Z(n7037) );
    GTECH_AND2 U2415 ( .A(n7009), .B(n7010), .Z(n7038) );
    GTECH_NAND2 U2416 ( .A(n7007), .B(n7008), .Z(n7035) );
    GTECH_AND2 U2417 ( .A(n7005), .B(n7006), .Z(n7036) );
    GTECH_AND2 U2418 ( .A(n7003), .B(n7004), .Z(n7033) );
    GTECH_AND2 U2419 ( .A(n7001), .B(n7002), .Z(n7034) );
    GTECH_AND2 U2420 ( .A(n7080), .B(n7079), .Z(n7095) );
    GTECH_AND2 U2421 ( .A(n7077), .B(n7078), .Z(n7096) );
    GTECH_NAND2 U2422 ( .A(n7076), .B(n7075), .Z(n7093) );
    GTECH_AND2 U2423 ( .A(n7073), .B(n7074), .Z(n7094) );
    GTECH_NAND2 U2424 ( .A(n7072), .B(n7071), .Z(n7091) );
    GTECH_AND2 U2425 ( .A(n7069), .B(n7070), .Z(n7092) );
    GTECH_NAND2 U2426 ( .A(n7068), .B(n7067), .Z(n7089) );
    GTECH_AND2 U2427 ( .A(n7065), .B(n7066), .Z(n7090) );
    GTECH_NAND2 U2428 ( .A(n7064), .B(n7063), .Z(n7087) );
    GTECH_AND2 U2429 ( .A(n7061), .B(n7062), .Z(n7088) );
    GTECH_NAND2 U2430 ( .A(n7060), .B(n7059), .Z(n7085) );
    GTECH_AND2 U2431 ( .A(n7057), .B(n7058), .Z(n7086) );
    GTECH_NAND2 U2432 ( .A(n7056), .B(n7055), .Z(n7083) );
    GTECH_AND2 U2433 ( .A(n7053), .B(n7054), .Z(n7084) );
    GTECH_AND2 U2434 ( .A(n7051), .B(n7052), .Z(n7081) );
    GTECH_AND2 U2435 ( .A(n7049), .B(n7050), .Z(n7082) );
    GTECH_AND2 U2436 ( .A(n7128), .B(n7127), .Z(n7143) );
    GTECH_AND2 U2437 ( .A(n7125), .B(n7126), .Z(n7144) );
    GTECH_AND2 U2438 ( .A(n7124), .B(n7123), .Z(n7141) );
    GTECH_AND2 U2439 ( .A(n7121), .B(n7122), .Z(n7142) );
    GTECH_NAND2 U2440 ( .A(n7120), .B(n7119), .Z(n7139) );
    GTECH_AND2 U2441 ( .A(n7117), .B(n7118), .Z(n7140) );
    GTECH_NAND2 U2442 ( .A(n7116), .B(n7115), .Z(n7137) );
    GTECH_AND2 U2443 ( .A(n7113), .B(n7114), .Z(n7138) );
    GTECH_NAND2 U2444 ( .A(n7112), .B(n7111), .Z(n7135) );
    GTECH_AND2 U2445 ( .A(n7109), .B(n7110), .Z(n7136) );
    GTECH_NAND2 U2446 ( .A(n7108), .B(n7107), .Z(n7133) );
    GTECH_AND2 U2447 ( .A(n7105), .B(n7106), .Z(n7134) );
    GTECH_NAND2 U2448 ( .A(n7103), .B(n7104), .Z(n7131) );
    GTECH_AND2 U2449 ( .A(n7102), .B(n7101), .Z(n7132) );
    GTECH_AND2 U2450 ( .A(n7100), .B(n7099), .Z(n7129) );
    GTECH_AND2 U2451 ( .A(n7097), .B(n7098), .Z(n7130) );
    GTECH_NOT U2452 ( .A(n6753), .Z(n6759) );
    GTECH_NAND2 U2453 ( .A(n6604), .B(\Exception_Index[3] ), .Z(n6482) );
    GTECH_AOI21 U2454 ( .A(n6519), .B(\Variables[0][-8][3]_wire ), .C(n6492), 
        .Z(n7156) );
    GTECH_AOI21 U2455 ( .A(n6519), .B(\Variables[0][-7][3]_wire ), .C(n6502), 
        .Z(n7151) );
    GTECH_AOI21 U2456 ( .A(n6519), .B(\Variables[0][-3][3]_wire ), .C(n6510), 
        .Z(n7153) );
    GTECH_NAND8 U2457 ( .A(n7172), .B(n7169), .C(n7166), .D(n7163), .E(n7160), 
        .F(n7157), .G(n7154), .H(n7150), .Z(n7192) );
    GTECH_NAND8 U2458 ( .A(n7189), .B(n7188), .C(n7187), .D(n7186), .E(n7185), 
        .F(n7184), .G(n7183), .H(n7181), .Z(n7194) );
    GTECH_AND_NOT U2459 ( .A(n6631), .B(n7319), .Z(n6643) );
    GTECH_AOI21 U2460 ( .A(n6336), .B(\Lower[0] ), .C(n6614), .Z(n6646) );
    GTECH_OR_NOT U2461 ( .A(\Upper[0] ), .B(n6336), .Z(n6645) );
    GTECH_AO21 U2462 ( .A(n6608), .B(n6607), .C(n6815), .Z(n6609) );
    GTECH_AO21 U2463 ( .A(n6813), .B(n6613), .C(n6814), .Z(n7324) );
    GTECH_AOI21 U2464 ( .A(n6816), .B(n7324), .C(n6817), .Z(n7325) );
    GTECH_OAI21 U2465 ( .A(n7325), .B(n6631), .C(n7326), .Z(n6617) );
    GTECH_NAND2 U2466 ( .A(n7176), .B(n7175), .Z(n7191) );
    GTECH_AO21 U2467 ( .A(n7193), .B(n7190), .C(n6825), .Z(n6441) );
    GTECH_AOI21 U2468 ( .A(n6519), .B(\Variables[0][-8][2]_wire ), .C(n6496), 
        .Z(n7202) );
    GTECH_AOI21 U2469 ( .A(n6519), .B(\Variables[0][-7][2]_wire ), .C(n6504), 
        .Z(n7197) );
    GTECH_AOI21 U2470 ( .A(n6519), .B(\Variables[0][-3][2]_wire ), .C(n6514), 
        .Z(n7198) );
    GTECH_NAND8 U2471 ( .A(n7218), .B(n7215), .C(n7212), .D(n7209), .E(n7206), 
        .F(n7203), .G(n7199), .H(n7196), .Z(n7235) );
    GTECH_NAND8 U2472 ( .A(n7232), .B(n7231), .C(n7230), .D(n7229), .E(n7228), 
        .F(n7227), .G(n7225), .H(n7223), .Z(n7237) );
    GTECH_OAI21 U2473 ( .A(n7327), .B(n6816), .C(n7328), .Z(n6620) );
    GTECH_NAND2 U2474 ( .A(n7222), .B(n7221), .Z(n7234) );
    GTECH_AO21 U2475 ( .A(n7236), .B(n7233), .C(n6825), .Z(n6443) );
    GTECH_AOI21 U2476 ( .A(n6519), .B(\Variables[0][-8][1]_wire ), .C(n6498), 
        .Z(n7242) );
    GTECH_AO21 U2477 ( .A(n6519), .B(\Variables[0][-7][1]_wire ), .C(n6506), 
        .Z(n7239) );
    GTECH_AOI21 U2478 ( .A(n6519), .B(\Variables[0][-3][1]_wire ), .C(n6516), 
        .Z(n7240) );
    GTECH_NAND8 U2479 ( .A(n7259), .B(n7256), .C(n7253), .D(n7250), .E(n7247), 
        .F(n7244), .G(n7241), .H(n7238), .Z(n7274) );
    GTECH_NAND8 U2480 ( .A(n7271), .B(n7270), .C(n7269), .D(n7268), .E(n7267), 
        .F(n7266), .G(n7265), .H(n7264), .Z(n7276) );
    GTECH_OAI21 U2481 ( .A(n6624), .B(n6813), .C(n7329), .Z(n6622) );
    GTECH_NAND2 U2482 ( .A(n7263), .B(n7262), .Z(n7273) );
    GTECH_AO21 U2483 ( .A(n7275), .B(n7272), .C(n6825), .Z(n6445) );
    GTECH_AOI21 U2484 ( .A(n6519), .B(\Variables[0][-8][0]_wire ), .C(n6500), 
        .Z(n7282) );
    GTECH_AOI21 U2485 ( .A(n6519), .B(\Variables[0][-7][0]_wire ), .C(n6508), 
        .Z(n7279) );
    GTECH_AOI21 U2486 ( .A(n6519), .B(\Variables[0][-3][0]_wire ), .C(n6518), 
        .Z(n7278) );
    GTECH_NAND8 U2487 ( .A(n7298), .B(n7295), .C(n7292), .D(n7289), .E(n7286), 
        .F(n7283), .G(n7280), .H(n7277), .Z(n7313) );
    GTECH_NAND8 U2488 ( .A(n7310), .B(n7309), .C(n7308), .D(n7307), .E(n7306), 
        .F(n7305), .G(n7304), .H(n7303), .Z(n7315) );
    GTECH_NAND2 U2489 ( .A(n7302), .B(n7301), .Z(n7312) );
    GTECH_AO21 U2490 ( .A(n7314), .B(n7311), .C(n6825), .Z(n6447) );
    GTECH_NAND3 U2491 ( .A(\NextInstruction[INSTRUCTION][3] ), .B(
        \NextInstruction[PARAMETER][3] ), .C(\NextInstruction[PARAMETER][2] ), 
        .Z(n7316) );
    GTECH_OAI21 U2492 ( .A(n6460), .B(n6664), .C(n6669), .Z(n7317) );
    GTECH_NAND3 U2493 ( .A(n6455), .B(n6453), .C(n6456), .Z(n6634) );
    GTECH_NAND5 U2494 ( .A(n6453), .B(n6450), .C(n6455), .D(n6615), .E(
        \NextInstruction[PARAMETER][1] ), .Z(n6632) );
    GTECH_OAI21 U2495 ( .A(n6448), .B(n6449), .C(n6430), .Z(n6636) );
    GTECH_XNOR3 U2496 ( .A(n6815), .B(n6608), .C(n6607), .Z(n6623) );
    GTECH_MUXI2 U2497 ( .A(n7319), .B(n6643), .S(n7325), .Z(n7326) );
    GTECH_MUX2 U2498 ( .A(\NextInstruction[INSTRUCTION][1] ), .B(n6627), .S(
        \NextInstruction[INSTRUCTION][3] ), .Z(n7180) );
    GTECH_MUXI2 U2499 ( .A(n6817), .B(n6611), .S(n7327), .Z(n7328) );
    GTECH_MUXI2 U2500 ( .A(n6814), .B(n6607), .S(n6624), .Z(n7329) );
    GTECH_OR3 U2501 ( .A(n6490), .B(\NextInstruction[INSTRUCTION][3] ), .C(
        n6660), .Z(n6846) );
    GTECH_NOT U2502 ( .A(n6662), .Z(n7178) );
    GTECH_NOT U2503 ( .A(RegularRegisterWrite), .Z(n6423) );
    GTECH_NOT U2504 ( .A(n6403), .Z(n6524) );
    GTECH_NOT U2505 ( .A(n6406), .Z(n6527) );
    GTECH_NOT U2506 ( .A(n6407), .Z(n6528) );
    GTECH_NOT U2507 ( .A(n6408), .Z(n6529) );
    GTECH_NOT U2508 ( .A(n6409), .Z(n6530) );
    GTECH_NOT U2509 ( .A(n6410), .Z(n6531) );
    GTECH_NOT U2510 ( .A(n6411), .Z(n6532) );
    GTECH_NOT U2511 ( .A(n6412), .Z(n6533) );
    GTECH_NOT U2512 ( .A(n6413), .Z(n6534) );
    GTECH_NOT U2513 ( .A(n6414), .Z(n6537) );
    GTECH_NOT U2514 ( .A(n6415), .Z(n6538) );
    GTECH_NOT U2515 ( .A(n6416), .Z(n6539) );
    GTECH_NOT U2516 ( .A(n6329), .Z(n6428) );
    GTECH_NOT U2517 ( .A(Write_wire), .Z(n6317) );
    GTECH_NOT U2518 ( .A(\RegularWriteRegister_Index[2] ), .Z(n6686) );
    GTECH_NOT U2519 ( .A(n6681), .Z(n6680) );
    GTECH_NOT U2520 ( .A(n6679), .Z(n7321) );
    GTECH_NOT U2521 ( .A(n6684), .Z(n7322) );
    GTECH_NOT U2522 ( .A(n6695), .Z(n7323) );
    GTECH_NOT U2523 ( .A(n6523), .Z(n6346) );
    GTECH_NOT U2524 ( .A(\Upper[0] ), .Z(n6785) );
    GTECH_NOT U2525 ( .A(n7145), .Z(n6996) );
    GTECH_NOT U2526 ( .A(n7147), .Z(n7045) );
    GTECH_NOT U2527 ( .A(n6775), .Z(n7146) );
    GTECH_NOT U2528 ( .A(n7151), .Z(n7182) );
    GTECH_NOT U2529 ( .A(n6820), .Z(n7224) );
    GTECH_NOT U2530 ( .A(n6784), .Z(n6789) );
    GTECH_NOT U2531 ( .A(n6795), .Z(n7201) );
    GTECH_NOT U2532 ( .A(n6788), .Z(n7152) );
    GTECH_NOT U2533 ( .A(n6747), .Z(n6997) );
    GTECH_NOT U2534 ( .A(\IPRELOAD_Table3551[2] ), .Z(n7149) );
    GTECH_NOT U2535 ( .A(n6604), .Z(n6318) );
    GTECH_NOT U2536 ( .A(Reset), .Z(n6472) );
    GTECH_NOT U2537 ( .A(n6605), .Z(n7148) );
    GTECH_NOT U2538 ( .A(n6613), .Z(n6624) );
    GTECH_NOT U2539 ( .A(n7324), .Z(n7327) );
    GTECH_NOT U2540 ( .A(n6330), .Z(n7226) );
    GTECH_NOT U2541 ( .A(n6435), .Z(n6439) );
    GTECH_NOT U2542 ( .A(\IRQ[0] ), .Z(n6325) );
    GTECH_FD1 \ClockCycleCount_reg[3]  ( .D(n7348), .CP(\CycleWaveform[5] ), 
        .QN(net108) );
    GTECH_FD1 \ClockCycleCount_reg[4]  ( .D(n7348), .CP(\CycleWaveform[5] ), 
        .QN(net109) );
    GTECH_FD1 \ClockCycleCount_reg[5]  ( .D(n7348), .CP(\CycleWaveform[5] ), 
        .QN(net110) );
    GTECH_FD1 \ClockCycleCount_reg[6]  ( .D(n7348), .CP(\CycleWaveform[5] ), 
        .QN(net111) );
    GTECH_FD1 \ClockCycleCount_reg[7]  ( .D(n7348), .CP(\CycleWaveform[5] ), 
        .QN(net112) );
    GTECH_FD1 \CycleWaveform_reg[5]  ( .D(\CycleWaveform34[5] ), .CP(
        InstructionReady), .Q(\CycleWaveform[5] ), .QN(n7330) );
    GTECH_FD1 \CycleWaveform_reg[4]  ( .D(\CycleWaveform34[4] ), .CP(
        InstructionReady), .Q(\CycleWaveform[4] ), .QN(n7331) );
    GTECH_FD1 \CycleWaveform_reg[3]  ( .D(\CycleWaveform34[3] ), .CP(
        InstructionReady), .Q(\CycleWaveform[3] ), .QN(n7332) );
    GTECH_FD1 \CycleWaveform_reg[2]  ( .D(\CycleWaveform34[2] ), .CP(
        InstructionReady), .Q(\CycleWaveform[2] ), .QN(n7333) );
    GTECH_FD1 \CycleWaveform_reg[1]  ( .D(\CycleWaveform34[1] ), .CP(
        InstructionReady), .Q(\CycleWaveform[1] ), .QN(n7334) );
    GTECH_FD1 \CycleWaveform_reg[0]  ( .D(\CycleWaveform34[0] ), .CP(
        InstructionReady), .QN(n7335) );
    GTECH_FD1S \ClockCycleCount_reg[0]  ( .D(ResetStarted), .TI(n7349), .TE(
        \sum1105[0] ), .CP(\CycleWaveform[5] ), .Q(\add_138/carry[1] ), .QN(
        n_399) );
    GTECH_FD1 \ClockCycleCount_reg[1]  ( .D(\ClockCycleCount621[1] ), .CP(
        \CycleWaveform[5] ), .Q(\ClockCycleCount[1] ), .QN(n_398) );
    GTECH_FD1 \ClockCycleCount_reg[2]  ( .D(\ClockCycleCount621[2] ), .CP(
        \CycleWaveform[5] ), .Q(\ClockCycleCount[2] ), .QN(n_397) );
    GTECH_FJK1S \TableSelect_reg[0]  ( .J(n7348), .K(n7348), .TI(
        \TableSelect667[0] ), .TE(\n668[3] ), .CP(\CycleWaveform[5] ), .Q(
        \TableSelect[0] ) );
    GTECH_FJK1S \TableSelect_reg[1]  ( .J(n7348), .K(n7348), .TI(
        \TableSelect667[1] ), .TE(\n668[3] ), .CP(\CycleWaveform[5] ), .Q(
        \TableSelect[1] ) );
    GTECH_FJK1S \TableSelect_reg[2]  ( .J(n7348), .K(n7348), .TI(
        \TableSelect667[2] ), .TE(\n668[3] ), .CP(\CycleWaveform[5] ), .Q(
        \gt_236/AEQB[2] ) );
    GTECH_FJK1S \TableSelect_reg[3]  ( .J(n7348), .K(n7348), .TI(
        \TableSelect667[3] ), .TE(\n668[3] ), .CP(\CycleWaveform[5] ), .Q(
        \TableSelect[3] ) );
    GTECH_FJK1S \RegularWriteRegister_Index_reg[0]  ( .J(n7348), .K(n7348), 
        .TI(\RegularWriteRegister_Index848[0] ), .TE(\n696[3] ), .CP(
        \CycleWaveform[5] ), .Q(\RegularWriteRegister_Index[0] ) );
    GTECH_FJK1S \RegularWriteRegister_Index_reg[1]  ( .J(n7348), .K(n7348), 
        .TI(\RegularWriteRegister_Index848[1] ), .TE(\n696[3] ), .CP(
        \CycleWaveform[5] ), .Q(\RegularWriteRegister_Index[1] ) );
    GTECH_FJK1S \RegularWriteRegister_Index_reg[2]  ( .J(n7348), .K(n7348), 
        .TI(\RegularWriteRegister_Index848[2] ), .TE(\n696[3] ), .CP(
        \CycleWaveform[5] ), .Q(\RegularWriteRegister_Index[2] ) );
    GTECH_FJK1S \RegularWriteRegister_Index_reg[3]  ( .J(n7348), .K(n7348), 
        .TI(\RegularWriteRegister_Index848[3] ), .TE(\n696[3] ), .CP(
        \CycleWaveform[5] ), .Q(\RegularWriteRegister_Index[3] ) );
    GTECH_FJK1S \Interrupt_Index_reg[0]  ( .J(n7348), .K(n7348), .TI(
        \NextInstruction[PARAMETER][0] ), .TE(\n706[3] ), .CP(
        \CycleWaveform[5] ), .Q(\Interrupt_Index[0] ) );
    GTECH_FJK1S \Interrupt_Index_reg[1]  ( .J(n7348), .K(n7348), .TI(
        \NextInstruction[PARAMETER][1] ), .TE(\n706[3] ), .CP(
        \CycleWaveform[5] ), .QN(n7336) );
    GTECH_FJK1S \Interrupt_Index_reg[2]  ( .J(n7348), .K(n7348), .TI(
        \NextInstruction[PARAMETER][2] ), .TE(\n706[3] ), .CP(
        \CycleWaveform[5] ), .Q(\Interrupt_Index[2] ) );
    GTECH_FJK1S \Interrupt_Index_reg[3]  ( .J(n7348), .K(n7348), .TI(
        \NextInstruction[PARAMETER][3] ), .TE(\n706[3] ), .CP(
        \CycleWaveform[5] ), .QN(n7337) );
    GTECH_FJK1S \Exception_Index_reg[0]  ( .J(n7348), .K(n7348), .TI(n7348), 
        .TE(n_358), .CP(\CycleWaveform[3] ), .Q(\Exception_Index[0] ) );
    GTECH_FJK1S \Exception_Index_reg[1]  ( .J(n7348), .K(n7348), .TI(n_324), 
        .TE(n_358), .CP(\CycleWaveform[3] ), .QN(n7338) );
    GTECH_FJK1S \Exception_Index_reg[2]  ( .J(n7348), .K(n7348), .TI(n_323), 
        .TE(n_358), .CP(\CycleWaveform[3] ), .Q(\Exception_Index[2] ) );
    GTECH_FJK1S \Exception_Index_reg[3]  ( .J(n7348), .K(n7348), .TI(n7348), 
        .TE(n_358), .CP(\CycleWaveform[3] ), .Q(\Exception_Index[3] ) );
    GTECH_FJK1S \IRQ_Index_reg[0]  ( .J(n7348), .K(n7348), .TI(n7348), .TE(
        n_726), .CP(\CycleWaveform[3] ), .Q(\IRQ_Index[0] ) );
    GTECH_FJK1S \IRQ_Index_reg[1]  ( .J(n7348), .K(n7348), .TI(n_566), .TE(
        n_726), .CP(\CycleWaveform[3] ), .QN(n7339) );
    GTECH_FJK1S \IRQ_Index_reg[2]  ( .J(n7348), .K(n7348), .TI(n_565), .TE(
        n_726), .CP(\CycleWaveform[3] ), .Q(\IRQ_Index[2] ) );
    GTECH_FJK1S \IRQ_Index_reg[3]  ( .J(n7348), .K(n7348), .TI(n_564), .TE(
        n_726), .CP(\CycleWaveform[3] ), .QN(n7340) );
    GTECH_FJK1S \IPRELOAD_Index_reg[0]  ( .J(n7348), .K(n7348), .TI(
        \IPRELOAD_Index3559[0] ), .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(
        \add_417/carry[1] ) );
    GTECH_FJK1S \IPRELOAD_Index_reg[1]  ( .J(n7348), .K(n7348), .TI(
        \IPRELOAD_Index3559[1] ), .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(
        \IPRELOAD_Index[1] ) );
    GTECH_FJK1S \IPRELOAD_Index_reg[2]  ( .J(n7348), .K(n7348), .TI(
        \IPRELOAD_Index3559[2] ), .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(
        \IPRELOAD_Index[2] ) );
    GTECH_FJK1S \IPRELOAD_Index_reg[3]  ( .J(n7348), .K(n7348), .TI(
        \IPRELOAD_Index3559[3] ), .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(
        \IPRELOAD_Index[3] ) );
    GTECH_FJK1S \MemoryPtr_reg[0]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[0] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[0] ) );
    GTECH_FJK1S \MemoryPtr_reg[1]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[1] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[1] ) );
    GTECH_FJK1S \MemoryPtr_reg[2]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[2] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[2] ) );
    GTECH_FJK1S \MemoryPtr_reg[3]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[3] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[3] ) );
    GTECH_FJK1S \MemoryPtr_reg[4]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[4] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[4] ) );
    GTECH_FJK1S \MemoryPtr_reg[5]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[5] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[5] ) );
    GTECH_FJK1S \MemoryPtr_reg[6]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[6] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[6] ) );
    GTECH_FJK1S \MemoryPtr_reg[7]  ( .J(n7348), .K(n7348), .TI(
        \MemoryPtr3672[7] ), .TE(\n3651[7] ), .CP(\CycleWaveform[2] ), .Q(
        \MemoryPtr[7] ) );
    GTECH_FJK1S \InstructionPtr_reg[0]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[0] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[0] ) );
    GTECH_FJK1S \InstructionPtr_reg[1]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[1] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[1] ) );
    GTECH_FJK1S \InstructionPtr_reg[2]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[2] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[2] ) );
    GTECH_FJK1S \InstructionPtr_reg[3]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[3] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[3] ) );
    GTECH_FJK1S \InstructionPtr_reg[4]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[4] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[4] ) );
    GTECH_FJK1S \InstructionPtr_reg[5]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[5] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[5] ) );
    GTECH_FJK1S \InstructionPtr_reg[6]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[6] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[6] ) );
    GTECH_FJK1S \InstructionPtr_reg[7]  ( .J(n7348), .K(n7348), .TI(
        \InstructionPtr3995[7] ), .TE(\n3996[7] ), .CP(\CycleWaveform[1] ), 
        .Q(\InstructionPtr[7] ) );
    GTECH_FJK1S Write_reg ( .J(n7348), .K(n7348), .TI(Write657), .TE(n658), 
        .CP(\CycleWaveform[5] ), .Q(Write_wire) );
    GTECH_FJK1S \Variables_reg[3][-6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-8][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-8][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-8][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-7][1] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-3][3] ), .TE(\n2831[0][-3][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][0][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][0][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][0][3]_wire ) );
    GTECH_FJK1S MemWait_reg ( .J(n7348), .K(n7348), .TI(\n3651[7] ), .TE(n3641
        ), .CP(\CycleWaveform[2] ), .QN(n7341) );
    GTECH_FJK1S \Variables_reg[0][6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-8][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-8][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-8][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-8][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-8][2] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-8][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-4][2]_wire ) );
    GTECH_FJK1S \IPRELOAD_Table_reg[1]  ( .J(n7348), .K(n7348), .TI(
        \IPRELOAD_Table3551[1] ), .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(
        \IPRELOAD_Table[1] ) );
    GTECH_FJK1S \Variables_reg[4][7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][0][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][0][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][0][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][0][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][0][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][0][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-5][2]_wire ) );
    GTECH_FJK1S Read_reg ( .J(n7348), .K(n7348), .TI(Read648), .TE(n658), .CP(
        \CycleWaveform[5] ), .Q(Read_wire) );
    GTECH_FJK1S \Variables_reg[1][-1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-8][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-8][0] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-8][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-8][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-8][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-8][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-7][3] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-8][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-8][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-8][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-3][1] ), .TE(\n2831[0][-3][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][0][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][0][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][0][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-3][0]_wire ) );
    GTECH_FJK1S IRQEnable_reg ( .J(n7348), .K(n7348), .TI(IRQEnable685), .TE(
        n686), .CP(\CycleWaveform[5] ), .Q(IRQEnable) );
    GTECH_FJK1S IRQJump_reg ( .J(n7348), .K(n7348), .TI(n_660), .TE(n7345), 
        .CP(\CycleWaveform[3] ), .Q(IRQJump) );
    GTECH_FJK1S \Variables_reg[1][2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][0][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][0][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][0][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-1][3]_wire ) );
    GTECH_FJK1 Condition_reg ( .J(n_4166), .K(n7348), .CP(\CycleWaveform[2] ), 
        .Q(Condition) );
    GTECH_FJK1S \Variables_reg[2][-2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-2][0]_wire ) );
    GTECH_FJK1S \Answer_reg[2]  ( .J(n7348), .K(n7348), .TI(\Answer639[2] ), 
        .TE(\n640[3] ), .CP(\CycleWaveform[5] ), .Q(\Lower[2] ) );
    GTECH_FJK1S \Variables_reg[2][-6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][7][1]_wire ) );
    GTECH_FD1S RegularJump_reg ( .D(n7348), .TI(n7345), .TE(
        \*cell*469/U11/Z_0 ), .CP(\CycleWaveform[5] ), .Q(RegularJump) );
    GTECH_FJK1S \Variables_reg[1][-6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][0][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][0][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][0][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][7][2]_wire ) );
    GTECH_FJK1S IRQReturnRegisterWrite_reg ( .J(n7348), .K(n7348), .TI(n_660), 
        .TE(n7345), .CP(\CycleWaveform[3] ), .QN(n7342) );
    GTECH_FJK1S \Variables_reg[0][-4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-8][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-8][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-8][2]_wire ) );
    GTECH_FJK1S \IRQ_reg[1]  ( .J(n7348), .K(n7348), .TI(n7348), .TE(n_690), 
        .CP(\CycleWaveform[3] ), .Q(\IRQ[1] ) );
    GTECH_FJK1S \Variables_reg[1][0][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][0][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][0][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][3][0]_wire ) );
    GTECH_FD1S ReturnJump_reg ( .D(n7348), .TI(n7345), .TE(\*cell*469/U10/Z_0 
        ), .CP(\CycleWaveform[5] ), .Q(ReturnJump) );
    GTECH_FJK1S \Variables_reg[1][-8][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-8][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-8][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-1][3]_wire ) );
    GTECH_FJK1S \Answer2_reg[0]  ( .J(n7348), .K(n7348), .TI(\Answer2629[0] ), 
        .TE(\n630[3] ), .CP(\CycleWaveform[5] ), .Q(\Upper[0] ) );
    GTECH_FJK1S \Variables_reg[0][-5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-1][1]_wire ) );
    GTECH_FJK1S \Answer2_reg[2]  ( .J(n7348), .K(n7348), .TI(\Answer2629[2] ), 
        .TE(\n630[3] ), .CP(\CycleWaveform[5] ), .Q(\Upper[2] ) );
    GTECH_FJK1S \Variables_reg[3][6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][5][2]_wire ) );
    GTECH_FD1S RegularReturnRegisterWrite_reg ( .D(n7348), .TI(n7345), .TE(
        \*cell*469/U9/Z_0 ), .CP(\CycleWaveform[5] ), .QN(n7343) );
    GTECH_FJK1S \Variables_reg[1][-8][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-8][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-8][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-8][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-8][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-8][0]_wire ) );
    GTECH_FJK1S \IRQ_reg[3]  ( .J(n7348), .K(n7348), .TI(n7348), .TE(n_692), 
        .CP(\CycleWaveform[3] ), .Q(\IRQ[3] ) );
    GTECH_FJK1S \Variables_reg[3][3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][0][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][0][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][0][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][0][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][0][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][0][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][4][0]_wire ) );
    GTECH_FD1S OpCodeRegisterWrite_reg ( .D(n7348), .TI(n_452), .TE(
        \*cell*469/U144/Z_0 ), .CP(\CycleWaveform[3] ), .Q(OpCodeRegisterWrite
        ) );
    GTECH_FJK1S \Variables_reg[0][1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][0][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][0][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][0][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-2][2]_wire ) );
    GTECH_FJK1S \Answer_reg[0]  ( .J(n7348), .K(n7348), .TI(\Answer639[0] ), 
        .TE(\n640[3] ), .CP(\CycleWaveform[5] ), .Q(\Lower[0] ) );
    GTECH_FJK1S \Variables_reg[4][1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-7][3]_wire ) );
    GTECH_FD1S RegularRegisterWrite_reg ( .D(n7348), .TI(n7345), .TE(
        \*cell*469/U7/Z_0 ), .CP(\CycleWaveform[5] ), .Q(RegularRegisterWrite)
         );
    GTECH_FJK1S \Variables_reg[2][-7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][0][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][0][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][0][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][0][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][0][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][0][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][1][0]_wire ) );
    GTECH_FJK1S \Answer_reg[1]  ( .J(n7348), .K(n7348), .TI(\Answer639[1] ), 
        .TE(\n640[3] ), .CP(\CycleWaveform[5] ), .Q(\Lower[1] ) );
    GTECH_FJK1S \Variables_reg[3][-5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][2][0]_wire ) );
    GTECH_FJK1S \Answer2_reg[3]  ( .J(n7348), .K(n7348), .TI(\Answer2629[3] ), 
        .TE(\n630[3] ), .CP(\CycleWaveform[5] ), .Q(\Upper[3] ) );
    GTECH_FJK1S \Variables_reg[1][5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-8][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-8][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-8][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-8][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-8][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-8][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][0][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][0][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][0][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][3][3]_wire ) );
    GTECH_FJK1S \IRQ_reg[2]  ( .J(n7348), .K(n7348), .TI(n7348), .TE(n_691), 
        .CP(\CycleWaveform[3] ), .Q(\IRQ[2] ) );
    GTECH_FJK1S \Variables_reg[0][-4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-8][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-8][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-8][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][0][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][0][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][0][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][3][1]_wire ) );
    GTECH_FJK1S \IRQ_reg[0]  ( .J(n7348), .K(n7348), .TI(n7348), .TE(n_689), 
        .CP(\CycleWaveform[3] ), .Q(\IRQ[0] ) );
    GTECH_FJK1S ResetStarted_reg ( .J(n7348), .K(n7348), .TI(Reset), .TE(n_168
        ), .CP(InstructionReady), .Q(ResetStarted), .QN(n7345) );
    GTECH_FJK1S \Variables_reg[1][-8][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-8][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-8][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][2][2]_wire ) );
    GTECH_FJK1S \Answer2_reg[1]  ( .J(n7348), .K(n7348), .TI(\Answer2629[1] ), 
        .TE(\n630[3] ), .CP(\CycleWaveform[5] ), .Q(\Upper[1] ) );
    GTECH_FJK1S \Variables_reg[1][5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-5][1]_wire ) );
    GTECH_FJK1S IRQWait_reg ( .J(n7348), .K(n7348), .TI(IRQWait611), .TE(n612), 
        .CP(\CycleWaveform[5] ), .QN(n7344) );
    GTECH_FJK1S \Variables_reg[3][-1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][0][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][0][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][0][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][1][2]_wire ) );
    GTECH_FJK1S \Answer_reg[3]  ( .J(n7348), .K(n7348), .TI(\Answer639[3] ), 
        .TE(\n640[3] ), .CP(\CycleWaveform[5] ), .Q(\Lower[3] ) );
    GTECH_FJK1S \IRQ_reg[4]  ( .J(n7348), .K(n7348), .TI(\IRQ2736[4] ), .TE(
        n_693), .CP(\CycleWaveform[3] ), .Q(\IRQ[4] ) );
    GTECH_FJK1S \Variables_reg[1][-6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][0][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][0][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][0][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][6][3]_wire ) );
    GTECH_FD1 OutOfRangeException_reg ( .D(OutOfRangeException2645), .CP(
        \CycleWaveform[4] ), .Q(n_324) );
    GTECH_FJK1S \Variables_reg[0][1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-7][2] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][7][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-8][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-8][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-8][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-3][0] ), .TE(\n2831[0][-3][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][0][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][0][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][0][0]_wire ) );
    GTECH_FD1S InterruptJump_reg ( .D(n7348), .TI(n7345), .TE(
        \*cell*469/U12/Z_0 ), .CP(\CycleWaveform[5] ), .Q(InterruptJump) );
    GTECH_FJK1S \Variables_reg[3][-3][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-3][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-3][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-7][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-7][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-7][3]_wire ) );
    GTECH_FJK1S IRQInProcess_reg ( .J(n7348), .K(n7348), .TI(IRQInProcess602), 
        .TE(n603), .CP(\CycleWaveform[5] ), .Q(IRQInProcess), .QN(n_452) );
    GTECH_FJK1S \Variables_reg[0][-2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-6][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-6][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-6][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-2][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-2][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-2][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][0][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][0][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][0][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-5][3]_wire ) );
    GTECH_FD1S ExceptionJump_reg ( .D(n7348), .TI(n_452), .TE(
        \*cell*469/U144/Z_0 ), .CP(\CycleWaveform[3] ), .Q(ExceptionJump) );
    GTECH_FJK1S \Variables_reg[1][-1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-8][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-8][1] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-8][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-4][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-4][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-4][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][3][0]_wire ) );
    GTECH_FJK1S \IPRELOAD_Table_reg[2]  ( .J(n7348), .K(n7348), .TI(
        \IPRELOAD_Table3551[2] ), .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(
        \IPRELOAD_Table[2] ) );
    GTECH_FJK1S \Variables_reg[0][6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][1][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][1][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][1][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][5][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][5][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][5][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-8][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-8][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-8][0]_wire ) );
    GTECH_FD1S BadOpCode_reg ( .D(n7348), .TI(n7345), .TE(\*cell*469/U6/Z_0 ), 
        .CP(\CycleWaveform[5] ), .QN(n7346) );
    GTECH_FJK1S \Variables_reg[1][-4][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-4][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-4][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-8][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-8][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-8][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-8][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-8][3] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-8][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][3][2]_wire ) );
    GTECH_FJK1S \IPRELOAD_Table_reg[0]  ( .J(n7348), .K(n7348), .TI(n7348), 
        .TE(n_4166), .CP(\CycleWaveform[2] ), .Q(\IPRELOAD_Table[0] ) );
    GTECH_FJK1S \Variables_reg[2][5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][6][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][6][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][6][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][2][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][2][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][2][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-3][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-3][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][7][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][7][0]_wire ) );
    GTECH_FD1S ExceptionReturnRegisterWrite_reg ( .D(n7348), .TI(n_452), .TE(
        \*cell*469/U144/Z_0 ), .CP(\CycleWaveform[3] ), .QN(n7347) );
    GTECH_FJK1S \Variables_reg[1][-5][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-5][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-5][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][-1][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][-1][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][-1][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][3][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][3][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][3][0]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-1][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-1][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-1][2]_wire ) );
    GTECH_FJK1S \Variables_reg[2][0][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][0][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][0][1]_wire ) );
    GTECH_FJK1S \Variables_reg[4][6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[0][7][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][7][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][7][2]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[2][4][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][4][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][4][3]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[2][-5][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[2][-5][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[2][-5][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-2][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-2][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-2][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][2][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][2][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][2][0]_wire ) );
    GTECH_FJK1S \Variables_reg[3][1][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][1][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][1][1]_wire ) );
    GTECH_FJK1S \Variables_reg[1][6][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][6][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][6][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-6][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-6][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-6][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][5][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][5][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][5][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][-7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][-7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][-7][1]_wire ) );
    GTECH_FJK1S IRQCLKEnable_reg ( .J(n7348), .K(n7348), .TI(IRQCLKEnable676), 
        .TE(n677), .CP(\CycleWaveform[5] ), .Q(IRQCLKEnable) );
    GTECH_FJK1S \Variables_reg[0][-7][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-7][0] ), .TE(\n2831[0][-8][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-7][0]_wire ) );
    GTECH_FJK1S \Variables_reg[1][3][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][3][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][3][3]_wire ) );
    GTECH_FJK1S \Variables_reg[1][7][1]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[1][7][1] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[1][7][1]_wire ) );
    GTECH_FJK1S \Variables_reg[3][4][0]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][4][0] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][4][0]_wire ) );
    GTECH_FJK1S \Variables_reg[4][-8][3]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[4][-8][3] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[4][-8][3]_wire ) );
    GTECH_FJK1S \Variables_reg[3][0][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[3][0][2] ), .TE(\n2831[4][7][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[3][0][2]_wire ) );
    GTECH_FJK1S \Variables_reg[0][-3][2]  ( .J(n7348), .K(n7348), .TI(
        \Variables2830[0][-3][2] ), .TE(\n2831[0][-3][3] ), .CP(
        \CycleWaveform[2] ), .Q(\Variables[0][-3][2]_wire ) );
    Neuron_DW01_inc_8_0 r228 ( .A({\InstructionPtr[7] , \InstructionPtr[6] , 
        \InstructionPtr[5] , \InstructionPtr[4] , \InstructionPtr[3] , 
        \InstructionPtr[2] , \InstructionPtr[1] , \InstructionPtr[0] }), .SUM(
        {\sum2964[7] , \sum2964[6] , \sum2964[5] , \sum2964[4] , \sum2964[3] , 
        \sum2964[2] , \sum2964[1] , \sum2964[0] }) );
    Neuron_DW02_mult_4_4_0 \Neuron_ALU_191/mul_168  ( .A({\Lower[3] , 
        \Lower[2] , \Lower[1] , \Lower[0] }), .B({\Upper[3] , \Upper[2] , 
        \Upper[1] , \Upper[0] }), .TC(n7349), .PRODUCT({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, \product1846[5] , \product1846[4] , 
        \product1846[3] , \product1846[2] , SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4}) );
endmodule

