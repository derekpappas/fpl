module as_tb  ; 

parameter period  = 100 ; 
  as    #( period  )
   DUT  ( ); 

endmodule

