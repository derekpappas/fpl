//test type : module_declaration
//vparser rule name : 
//author : Codrin
(* a *)
(* a = 1 *)
module declaration_010;
endmodule
