//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : agent_long_reach.v
//FILE GENERATED ON : Thu Aug 14 15:17:29 2008

`include "defines.v"

module agent_long_reach();
// Location of source csl unit: file name = generated/agent_cl.csl line number = 72
  `include "agent_long_reach.logic.v"
endmodule

