`include "defines.v"

module u5();
// Location of source csl unit: file name = ar16.csl line number = 51
  `include "u5.logic.v"
endmodule

