//test type : module_or_generate_item ::= local_parameter_declaration
//vparser rule name : 
//author : Codrin
module test_0550;
 (* starts = "0" , waits = 5 *)
 localparam a = 8'b10101010, b = 1'hZ, c = 5;
endmodule
