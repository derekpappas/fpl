// Test type: disable_statement - disable hierarchical block id
// Vparser rule name:
// Author: andreib
module disable_statement2;

initial begin: TEST
disable TEST;
end
endmodule
