// Test type: Hex Numbers - signed value
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8'sh3F;
endmodule
