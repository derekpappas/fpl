// Test type: Real numbers - all numbers
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1234567890.1234567890e9;
endmodule
