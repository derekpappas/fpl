// Test type: seq_block - begin - 1 statement - end
// Vparser rule name:
// Author: andreib
module seq_block3;
reg a;
initial begin
	a=1'b1;
	end
endmodule
