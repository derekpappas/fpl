`include "defines.v"

module mem();
// Location of source csl unit: file name = parameter_test9.csl line number = 3
// The depth of memory module mem is of illegal type. Depth set to 1.
// The width of memory module mem is of illegal type. Width set to 1.
  parameter data_w = 4;
  parameter addr_w = 8;
  endmodule

