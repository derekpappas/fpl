--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : ssm.vh
--FILE GENERATED ON : Sat May  1 19:39:32 2010

Va2r_tap.vhd
arm.vhd
cmpr.vhd
dsp.vhd
dummy_unit_synth_removes.vhd
eu.vhd
h264.vhd
im.vhd
me.vhd
pc.vhd
rf.vhd
ssm.vhd
ssm_master.vhd
wb.vhd
