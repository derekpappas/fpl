`celldefine
module uid;
endmodule
`include "../legal/celldef08.v"
module sguid;
endmodule
`include "../legal/celldef07.v"
