`define operator =
module x;
reg a,b;
wire c;
if( a =`operator b);
endmodule
