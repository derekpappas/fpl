// Test type: nonblocking_assignment - expression
// Vparser rule name:
// Author: andreib
module nonblocking_assignment1;
reg a;
initial a<=1'b1;
endmodule
