`include "defines.v"

module a1(p1);
// Location of source csl unit: file name = f2a_p_out.csl line number = 3
  output [4 - 1:0] p1;
  `include "a1.logic.v"
endmodule

