`default_nettype none
`default_nettype trireg
module x;
`default_nettype none`resetall
