`define __ numero1
`define \_ _ `a(_)
`define a(_)\
this is a macro\
continued on the next line _\comment? \
a(_)
`a(\)
module x`__(y);
input y;
reg y;
endmodule //end of module xnumero1(y)

