u1.vhd
u2.vhd
