//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : eth_bridge.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module eth_bridge(eb_emdummy4,
                  lbdummy2);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 47
  input lbdummy2;
  output eb_emdummy4;
  `include "eth_bridge.logic.v"
endmodule

