// Test type: Continuous assignment - st1, st0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous331;
wire a;
assign (strong1, strong0) a=1'b1;
endmodule
