//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : i2c_lba.v
//FILE GENERATED ON : Thu Jun 19 15:32:42 2008

`include "defines.v"

module i2c_lba(lbdummy3,
               lbadummy2);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 29
  input lbadummy2;
  output lbdummy3;
  `include "i2c_lba.logic.v"
endmodule

