ua.vhd
ub.vhd
uc.vhd
ud.vhd
ue.vhd
ude.vhd
uf.vhd
ar15a.vhd
