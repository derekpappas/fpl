//this is a celldefine valid test
module mod;
`celldefine
wire x;
`resetall
endmodule
