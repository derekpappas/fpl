//THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
//COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
//OUTPUT FILE NAME  : nina.v
//FILE GENERATED ON : Tue Jun 17 01:23:46 2008

`include "defines.v"

module nina(lbadummy3);
// Location of source csl unit: file name = generated/msi_phase_1.csl line number = 42
  input lbadummy3;
  `include "nina.logic.v"
endmodule

