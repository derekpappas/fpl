-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./proc_ring_cslc_generated/code/vhdl/qm.vhd
-- FILE GENERATED ON : Wed Jul  9 20:26:20 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \qm\ is
  port(\dwaddr\ : in csl_bit_vector(17 downto 0);
       \dwdata\ : in csl_bit_vector(31 downto 0);
       \dwwr\ : out csl_bit);
begin
end entity;

architecture \qm_logic\ of \qm\ is
begin
end architecture;

