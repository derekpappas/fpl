`include "defines.v"

module b0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 7
  input [1 - 1:0] ar_sa0_s10;
  a0 a0(.sa0(ar_sa0_s10));
  `include "b0.logic.vh"
endmodule

