MAC_rx.vhd
MAC_tx.vhd
Phy_int.vhd
Reg_int.vhd
RMON.vhd
eth_miim.vhd
Clk_ctrl.vhd
MAC_top.vhd
