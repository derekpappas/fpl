// Test type: Octal Numbers - space between size and base
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=24 'o23454761;
endmodule
