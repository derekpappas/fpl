// Test type: Continuous assignment - wk1, h0 - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous601;
wire a;
assign (weak1, highz0) a=1'b1;
endmodule
