`include "defines.v"

module crc();
// Location of source csl unit: file name = IPX2400.csl line number = 50
  `include "crc.logic.v"
endmodule

