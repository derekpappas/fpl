// Test type: Octal Numbers - signed octal number
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=9'so123;
endmodule
