`include "defines.v"

module d1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 201
  output [1 - 1:0] ar_sa0_s10;
  c1 c10(.ar_sa0_s10(ar_sa0_s10));
  `include "d1.logic.vh"
endmodule

