// Dummy
// By Claudiu
// Used for compatibility issues

module lpm_decode;


endmodule
