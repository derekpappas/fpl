-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./msi_rx_cslc_generated/code/vhdl/ddr_buf_ctrl.vhd
-- FILE GENERATED ON : Thu Jun 19 15:32:42 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \ddr_buf_ctrl\ is
  port(\lbdummy3\ : out csl_bit;
       \lbadummy2\ : in csl_bit);
begin
end entity;

architecture \ddr_buf_ctrl_logic\ of \ddr_buf_ctrl\ is
begin
end architecture;

