//test type : number binary_operator_<= number
//vparser rule name : 
//author : Bogdan Mereghea
module binary_operator39;
    wire a;
    assign a = 1'b1 <= 1'b0;
endmodule
