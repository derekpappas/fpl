module testbench_charge_strength;
  charge_strength0 charge_strength_instance0();
  charge_strength0 charge_strength_instance1();
  charge_strength0 charge_strength_instance2();
  charge_strength0 charge_strength_instance3();
  charge_strength0 charge_strength_instance4();
  charge_strength0 charge_strength_instance5();
  charge_strength0 charge_strength_instance6();
  charge_strength0 charge_strength_instance7();
  charge_strength0 charge_strength_instance8();
  charge_strength0 charge_strength_instance9();
  charge_strength0 charge_strength_instance10();
  charge_strength0 charge_strength_instance11();
endmodule
//author : andreib
module charge_strength0;
trireg (small) a;
endmodule
//author : andreib
module charge_strength1;
trireg (small ) a;
endmodule
//author : andreib
module charge_strength2;
trireg ( small) a;
endmodule
//author : andreib
module charge_strength3;
trireg ( small ) a;
endmodule
//author : andreib
module charge_strength4;
trireg (medium) a;
endmodule
//author : andreib
module charge_strength5;
trireg (medium ) a;
endmodule
//author : andreib
module charge_strength6;
trireg ( medium) a;
endmodule
//author : andreib
module charge_strength7;
trireg ( medium ) a;
endmodule
//author : andreib
module charge_strength8;
trireg (large) a;
endmodule
//author : andreib
module charge_strength9;
trireg (large ) a;
endmodule
//author : andreib
module charge_strength10;
trireg ( large) a;
endmodule
//author : andreib
module charge_strength11;
trireg ( large ) a;
endmodule

