// Test type: net_assignment - binary operator, no attribute instance
// Vparser rule name:
// Author: andreib
module netasign5;
wire a,b,c;
assign a=b+c;
endmodule
