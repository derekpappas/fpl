module x;
`default_nettype
