// Dummy by Claudiu

module GTECH_ADD_AB;
endmodule

module GTECH_NOT;
endmodule

module GTECH_OAI2N2;
endmodule

module GTECH_ADD_ABC;
endmodule

module GTECH_AND2;
endmodule

module GTECH_AND_NOT;
endmodule

module GTECH_XOR3;
endmodule

module GTECH_NOR2;
endmodule

module GTECH_NAND2;
endmodule

module GTECH_ZERO;
endmodule

module GTECH_ONE;
endmodule

module GTECH_OR_NOT;
endmodule

module TECH_OR2;
endmodule

module GTECH_OAI21;
endmodule

module GTECH_AO21;
endmodule

module GTECH_0A21;
endmodule

module GTECH_AO22;
endmodule

module GTECH_OR2;
endmodule

module GTECH_OA21;
endmodule

module GTECH_OAI22;
endmodule

module GTECH_NAND3;
endmodule

module GTECH_OR3;
endmodule

module GTECH_NAND4;
endmodule

module GTECH_NOR3;
endmodule

module GTECH_AOI222;
endmodule

module GTECH_AND3;
endmodule

module GTECH_AND8;
endmodule

module GTECH_MAJ23;
endmodule

module GTECH_MUXI2;
endmodule

module TECH_AND4;
endmodule

module GTECH_AOI2N2;
endmodule

module GTECH_AND5;
endmodule

module GTECH_AOI21;
endmodule

module GTECH_AOI22;
endmodule

module GTECH_AND4;
endmodule

module GTECH_MUX2;
endmodule

module GTECH_OA22;
endmodule

module GTECH_NAND5;
endmodule

module GTECH_NAND8;
endmodule

module GTECH_XNOR3;
endmodule

module GTECH_FD1;
endmodule

module GTECH_FD1S;
endmodule

module GTECH_FJK1S;
endmodule

module GTECH_FJK1;
endmodule
