module testbench_function_declaration000;
    function_declaration001 function_declaration1_instance001();
endmodule

module function_declaration001;
reg a,b,c;
function automatic signed time function_identifier0123456789 ; 
input d; 
(* b , c *) (* b , c *) (* b , c *) input time port_identifier_abc , _port_identifier_ABC ; 
begin
a=1'b1;
a=a+1'b1;
end
 endfunction
endmodule
