// Test type: Real numbers - 1 number
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1.3;
endmodule
