`include "defines.v"

module dramctrl();
// Location of source csl unit: file name = IPX2400.csl line number = 95
  `include "dramctrl.logic.v"
endmodule

