module unit_b;
  wire sgn_in;
  reg sgn_out;
endmodule