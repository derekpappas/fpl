`include "defines.v"

module l1(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 250
  output [1 - 1:0] ar_sa0_s10;
  k1 k10(.ar_sa0_s10(ar_sa0_s10));
  `include "l1.logic.vh"
endmodule

