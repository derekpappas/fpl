// Test type: Decimal Numbers - lower case decimal base
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=5'd16;
endmodule
