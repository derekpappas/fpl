// Test type: initial statement - loop_statement - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon16;
reg [7:0]a;
initial forever a=2;
endmodule
