-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./b_cslc_generated/code/vhdl/b_a0.vhd
-- FILE GENERATED ON : Mon Feb 16 21:25:24 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \b_a0\ is
  port(\x\ : in csl_bit);
begin
end entity;

architecture \b_a0_logic\ of \b_a0\ is
begin
end architecture;

