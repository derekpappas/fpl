// Test type: Continuous assignment - list_of_net_assignments - 1 element
// Vparser rule name:
// Author: andreib
module continuous1;
wire a;
assign a=1'b1;
endmodule
