// Test type: Constant Expression - primary - param
// Vparser rule name:
// Author: andreib
module constantexpression;
parameter test=0;
endmodule
