// Test type: Binary Numbers - Underscore within value
// Vparser rule name: Numbers
// Author: andreib
module binary_num;
wire a;
assign a=6'b011_010_;
endmodule
