`include "defines.v"

module j0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 63
  input [1 - 1:0] ar_sa0_s10;
  i0 i0(.ar_sa0_s10(ar_sa0_s10));
  `include "j0.logic.vh"
endmodule

