-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./v_top_cslc_generated/code/vhdl/gpio.vhd
-- FILE GENERATED ON : Wed Sep 17 15:37:32 2008
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \gpio\ is
  port(\gp_in\ : out csl_bit;
       \gp_out\ : in csl_bit;
       \gp_en\ : in csl_bit);
begin
end entity;

architecture \gpio_logic\ of \gpio\ is
begin
end architecture;

