// Test type: initial statement - event_trigger - no attribute instance
// Vparser rule name:
// Author: andreib
module initcon13;
event a;
initial ->a;
endmodule
