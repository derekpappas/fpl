//this is a celldefine legal test
`celldefine
module mymodule;
endmodule

