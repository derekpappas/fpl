reg1.vhd
u1.vhd
