// Test type: Octal Numbers - underscores within octal value
// Vparser rule name: Numbers
// Author: andreib
module octal_num;
wire a;
assign a=9'o1_52_;
endmodule
