// Test type: loop statement - repeat
// Vparser rule name:
// Author: andreib
module loop_statement2;
reg a;
initial repeat(4) a=a+1;
endmodule
