//this is a celldefine legal test
module mod;
/**//***//**/`celldefine/***///sa
module mymodule;
endmodule
/****/`endcelldefine//haha
/*hihi*/endmodule
