//test type : specify_block_declaration
//author : Dramba Doru-Gabriel
module specify_block20(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; endspecify
endmodule
module specify_block21(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block22(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block23(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block24(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block25(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block26(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block27(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block28(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block29(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block210(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block211(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block212(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block213(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block214(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block215(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block216(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block217(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block218(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block219(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block220(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block221(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block222(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block223(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block224(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block225(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block226(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block227(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block228(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block229(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block230(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block231(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; endspecify
endmodule
module specify_block232(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block233(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block234(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block235(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block236(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block237(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block238(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block239(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block240(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block241(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block242(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block243(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block244(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block245(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block246(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block247(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block248(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block249(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block250(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block251(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block252(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block253(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block254(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block255(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block256(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block257(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block258(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block259(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block260(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block261(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block262(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block263(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block264(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block265(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block266(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block267(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block268(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block269(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block270(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block271(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block272(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block273(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block274(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block275(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block276(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block277(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block278(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block279(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block280(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block281(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block282(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block283(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block284(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block285(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block286(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block287(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block288(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block289(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block290(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block291(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block292(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block293(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block294(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block295(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block296(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block297(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block298(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block299(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2100(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2101(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2102(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2103(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2104(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2105(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2106(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2107(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2108(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2109(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2110(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2111(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2112(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2113(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2114(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2115(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2116(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2117(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2118(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2119(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2120(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2121(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2122(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2123(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2124(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2125(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2126(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2127(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2128(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2129(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2130(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2131(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2132(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2133(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2134(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2135(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2136(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2137(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2138(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2139(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2140(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2141(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2142(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2143(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2144(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2145(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2146(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2147(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2148(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2149(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2150(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2151(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2152(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2153(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2154(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2155(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2156(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2157(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2158(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2159(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2160(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2161(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2162(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2163(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2164(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2165(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2166(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2167(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2168(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2169(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2170(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2171(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2172(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2173(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2174(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2175(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2176(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2177(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2178(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2179(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2180(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2181(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2182(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2183(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2184(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2185(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam ter1 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2186(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2187(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2188(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2189(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2190(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2191(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2192(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2193(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2194(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2195(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2196(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2197(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2198(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2199(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2200(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2201(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2202(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2203(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2204(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2205(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2206(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2207(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2208(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2209(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2210(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2211(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2212(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2213(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2214(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2215(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2216(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2217(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; endspecify
endmodule
module specify_block2218(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2219(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2220(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2221(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2222(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2223(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2224(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2225(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2226(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2227(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2228(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2229(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2230(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2231(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2232(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2233(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2234(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2235(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2236(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2237(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2238(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2239(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2240(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2241(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2242(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2243(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2244(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2245(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2246(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2247(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2248(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2249(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2250(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2251(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2252(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2253(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2254(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2255(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2256(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2257(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2258(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2259(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2260(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2261(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2262(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2263(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2264(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2265(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2266(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2267(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2268(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2269(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2270(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2271(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2272(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2273(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2274(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2275(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2276(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2277(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2278(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2279(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2280(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2281(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2282(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2283(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2284(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2285(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2286(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2287(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2288(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2289(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2290(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2291(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2292(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2293(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2294(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2295(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2296(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2297(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2298(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2299(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2300(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2301(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2302(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2303(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2304(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2305(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2306(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2307(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2308(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2309(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2310(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2311(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2312(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2313(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2314(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2315(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2316(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2317(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2318(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2319(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2320(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2321(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2322(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2323(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2324(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2325(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2326(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2327(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2328(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2329(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2330(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2331(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2332(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2333(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2334(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2335(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2336(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2337(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2338(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2339(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2340(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2341(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2342(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2343(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2344(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2345(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2346(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2347(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2348(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2349(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2350(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2351(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2352(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2353(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2354(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2355(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2356(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2357(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2358(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2359(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2360(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2361(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2362(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2363(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2364(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2365(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2366(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2367(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2368(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2369(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2370(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2371(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2372(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2373(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2374(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2375(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2376(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2377(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2378(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2379(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2380(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2381(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2382(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2383(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2384(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2385(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2386(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2387(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2388(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2389(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2390(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2391(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2392(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2393(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2394(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2395(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2396(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2397(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2398(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2399(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2400(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2401(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2402(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2403(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; endspecify
endmodule
module specify_block2404(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2405(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2406(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2407(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2408(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2409(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2410(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2411(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2412(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2413(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2414(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2415(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2416(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2417(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2418(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2419(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2420(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2421(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2422(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2423(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2424(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2425(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2426(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2427(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2428(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2429(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2430(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2431(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2432(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2433(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2434(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2435(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2436(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2437(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2438(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2439(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2440(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2441(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2442(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2443(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2444(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2445(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2446(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2447(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2448(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2449(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2450(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2451(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2452(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2453(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2454(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2455(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2456(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2457(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2458(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2459(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2460(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2461(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2462(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2463(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2464(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2465(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2466(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2467(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2468(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2469(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2470(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2471(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2472(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2473(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2474(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2475(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2476(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2477(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2478(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2479(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2480(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2481(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2482(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2483(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2484(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2485(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2486(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2487(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2488(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2489(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2490(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2491(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2492(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2493(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2494(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2495(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2496(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2497(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2498(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2499(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2500(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2501(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2502(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2503(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2504(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2505(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2506(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2507(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2508(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2509(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2510(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2511(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2512(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2513(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2514(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2515(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2516(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2517(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2518(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2519(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2520(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2521(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2522(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2523(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2524(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2525(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2526(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2527(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2528(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2529(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2530(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2531(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2532(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2533(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2534(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2535(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2536(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2537(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2538(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2539(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2540(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2541(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2542(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2543(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2544(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2545(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2546(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2547(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2548(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2549(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2550(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2551(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2552(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2553(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2554(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2555(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2556(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2557(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2558(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2559(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2560(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2561(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2562(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2563(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2564(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2565(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2566(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2567(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2568(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2569(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2570(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2571(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2572(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2573(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2574(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2575(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2576(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2577(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2578(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2579(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2580(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2581(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2582(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2583(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2584(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2585(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2586(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2587(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2588(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2589(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; endspecify
endmodule
module specify_block2590(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2591(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2592(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2593(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2594(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2595(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2596(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2597(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2598(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2599(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2600(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2601(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2602(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2603(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2604(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2605(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2606(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2607(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2608(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2609(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2610(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2611(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2612(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2613(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2614(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2615(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2616(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2617(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2618(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2619(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2620(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2621(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2622(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2623(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2624(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2625(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2626(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2627(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2628(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2629(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2630(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2631(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2632(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2633(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2634(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2635(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2636(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2637(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2638(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2639(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2640(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2641(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2642(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2643(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2644(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2645(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2646(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2647(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2648(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2649(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2650(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2651(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2652(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2653(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2654(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2655(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2656(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2657(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2658(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2659(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2660(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2661(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2662(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2663(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2664(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2665(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2666(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2667(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2668(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2669(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2670(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2671(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2672(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2673(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2674(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2675(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2676(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2677(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2678(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2679(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2680(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2681(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2682(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2683(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2684(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2685(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2686(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2687(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2688(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2689(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2690(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2691(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2692(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2693(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2694(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2695(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2696(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2697(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2698(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2699(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2700(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2701(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2702(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2703(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2704(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2705(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2706(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2707(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2708(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2709(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2710(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2711(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2712(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2713(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2714(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2715(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2716(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2717(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2718(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2719(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2720(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2721(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2722(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2723(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2724(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2725(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2726(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2727(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2728(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2729(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2730(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2731(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2732(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2733(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2734(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2735(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2736(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2737(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2738(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2739(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2740(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2741(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2742(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2743(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2744(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2745(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2746(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2747(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2748(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2749(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2750(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2751(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2752(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2753(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2754(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2755(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2756(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2757(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2758(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2759(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2760(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2761(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2762(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2763(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2764(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2765(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2766(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2767(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2768(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2769(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2770(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2771(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2772(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2773(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2774(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2775(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; endspecify
endmodule
module specify_block2776(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2777(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2778(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2779(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2780(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2781(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2782(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2783(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2784(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2785(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2786(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2787(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2788(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2789(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2790(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2791(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2792(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2793(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2794(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2795(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2796(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2797(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2798(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2799(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2800(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2801(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2802(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2803(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2804(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2805(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter2 = 1 ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2806(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2807(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2808(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2809(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2810(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2811(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2812(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2813(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2814(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2815(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2816(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2817(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2818(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2819(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2820(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2821(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2822(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2823(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2824(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2825(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2826(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2827(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2828(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2829(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2830(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2831(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2832(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2833(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2834(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2835(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2836(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2837(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2838(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2839(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2840(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2841(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2842(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2843(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2844(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2845(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2846(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2847(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2848(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2849(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2850(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2851(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2852(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2853(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2854(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2855(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2856(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2857(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2858(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2859(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2860(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2861(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2862(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2863(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2864(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2865(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2866(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2867(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2868(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2869(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2870(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2871(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2872(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2873(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2874(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2875(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2876(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2877(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2878(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2879(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2880(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2881(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2882(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2883(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2884(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2885(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2886(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2887(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2888(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2889(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2890(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2891(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2892(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2893(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2894(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2895(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2896(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2897(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2898(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2899(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2900(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 ; endspecify
endmodule
module specify_block2901(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , ter4 = 1 ; endspecify
endmodule
module specify_block2902(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2903(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2904(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2905(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam ter3 = 1 , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2906(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2907(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2908(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2909(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2910(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2911(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2912(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2913(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2914(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2915(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2916(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2917(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2918(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2919(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2920(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2921(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2922(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2923(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2924(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
module specify_block2925(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , ter4 = 1 ; endspecify
endmodule
module specify_block2926(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 ) ; endspecify
endmodule
module specify_block2927(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$=( 10 , 10 ) ; endspecify
endmodule
module specify_block2928(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 ) ; endspecify
endmodule
module specify_block2929(inoutPortIdentifier,outputPortIdentifier,outputPortIdentifier2);
  inout inoutPortIdentifier;
  output outputPortIdentifier;
  output [14:0] outputPortIdentifier2;
  specify specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; specparam PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) , PATHPULSE$inoutPortIdentifier$outputPortIdentifier=( 10 , 10 ) ; endspecify
endmodule
