// Dummy
// By Claudiu
// Used for compatibility issues

module opndrn;


endmodule
