//test type : port_declaration
//vparser rule name : 
//author : Codrin
module declaration_090(x);
 (* a = 1, b *) input x;
endmodule
