`include "defines.v"

module im();
// Location of source csl unit: file name = /Volumes/s2/unfuddle_ssm_repo/ssm_ssmrepo/ssm/hw/ssm/ssm_demo.csl line number = 93
  `include "im.logic.vh"
endmodule

