module a(x);
output x;
endmodule
