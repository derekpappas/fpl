//test type : operator_^ system_funtion_call
//vparser rule name : 
//author : Bogdan Mereghea
module unary_operator64;
    wire a;
    assign a = ^$random;
endmodule
