// Test type: Real numbers - underscores within
// Vparser rule name: Numbers
// Author: andreib
module real_num;
wire a;
assign a=1234_567_.1_2_e1_23_;
endmodule
