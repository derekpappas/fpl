// Test type: Hex Numbers - space between size and base
// Vparser rule name: Numbers
// Author: andreib
module hex_num;
wire a;
assign a=8 'h78;
endmodule
