// Test type: Decimal Numbers - no size decimal base lower case
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a='d79;
endmodule
