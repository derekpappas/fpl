//test type : module_declaration
//vparser rule name : 
//author : Codrin
(* a *)
module declaration_000;
endmodule
