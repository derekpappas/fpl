-------------------------------------------------------------------------------
-- THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
-- COPYRIGHT (c) 2006-2008 FastpathLogic Inc
-- FILE NAME         : ./u_dep_cslc_generated/code/vhdl/u_ff.vhd
-- FILE GENERATED ON : Mon Feb 16 21:29:41 2009
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

library csl_util;
use csl_util.csl_util_package.all;

entity \u_ff\ is
  generic(\width\ : csl_integer := 10#1#);
  port(\d\ : in csl_bit_vector(\width\ - 10#1# downto 10#0#);
       \q\ : out csl_bit_vector(\width\ - 10#1# downto 10#0#);
       \reset\ : in csl_bit;
       \enable\ : in csl_bit;
       \clk\ : in csl_bit);
begin
end entity;

architecture \u_ff_logic\ of \u_ff\ is
begin
end architecture;

