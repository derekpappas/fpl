--THIS CODE WAS GENERATED USING THE FASTPATHLOGIC HDL COMPILER
--COPYRIGHT (c) 2006, 2007 FastpathLogic Inc
--OUTPUT FILE NAME  : eu.vhd
--FILE GENERATED ON : Sat May  1 19:39:32 2010


library ieee ; 
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all; 
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
 
use work.csl_util_package.all;

entity eu is 

-- Location of source csl unit: file name = /Volumes/s2/unfuddle_ssm_repo/ssm_ssmrepo/ssm/hw/ssm/ssm_demo.csl line number = 91
end eu ; 

 architecture  arch_eu of eu is 

dummy1_master_ifc_address : in   csl_bit_vector(0 downto 0);
dummy1_master_ifc_write_data : in   csl_bit_vector(0 downto 0);
dummy1_master_ifc_read : in   csl_bit_vector(0 downto 0);
dummy1_master_ifc_write : in   csl_bit_vector(0 downto 0);
dummy2_master_ifc_address : in   csl_bit_vector(0 downto 0);
dummy2_master_ifc_write_data : in   csl_bit_vector(0 downto 0);
dummy2_master_ifc_read : in   csl_bit_vector(0 downto 0);
dummy2_master_ifc_write : in   csl_bit_vector(0 downto 0);
dummy3_master_ifc_address : in   csl_bit_vector(0 downto 0);
dummy3_master_ifc_write_data : in   csl_bit_vector(0 downto 0);
dummy3_master_ifc_read : in   csl_bit_vector(0 downto 0);
dummy3_master_ifc_write : in   csl_bit_vector(0 downto 0);
dummy1_master_ifc_read_data : out   csl_bit_vector(0 downto 0);
dummy1_master_ifc_ready : out   csl_bit_vector(0 downto 0);
dummy1_master_ifc_error : out   csl_bit_vector(0 downto 0);
dummy2_master_ifc_read_data : out   csl_bit_vector(0 downto 0);
dummy2_master_ifc_ready : out   csl_bit_vector(0 downto 0);
dummy2_master_ifc_error : out   csl_bit_vector(0 downto 0);
dummy3_master_ifc_read_data : out   csl_bit_vector(0 downto 0);
dummy3_master_ifc_ready : out   csl_bit_vector(0 downto 0);
dummy3_master_ifc_error : out   csl_bit_vector(0 downto 0) 
 begin 

 end  arch_eu ; 
