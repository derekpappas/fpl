`include "defines.v"

module o0(ar_sa0_s10);
// Location of source csl unit: file name = temp.csl line number = 101
  input [1 - 1:0] ar_sa0_s10;
  n0 n0(.ar_sa0_s10(ar_sa0_s10));
  `include "o0.logic.vh"
endmodule

