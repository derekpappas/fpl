//test type : non_port_module_item ::= parameter_declaration
//vparser rule name : 
//author : Codrin
module test_0380;
 (* debug = 1, test *)
 parameter msb = 7;
endmodule
