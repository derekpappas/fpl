// Test type: Decimal Numbers - Simple decimal number
// Vparser rule name: Numbers
// Author: andreib
module decimal_num;
wire a;
assign a=2;
endmodule
